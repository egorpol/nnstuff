BZh91AY&SY��{0*_�ryg��������� @ b!>� 
� �( ��H P  ��%@J %ATB%R
@ R@  �����*��EP$HUH  
RIE%!B���UQATD( 

��
�@�D�";��� P��P���I(
)@   HQT��(��*�) ���
 �
�%{�%*�{��`�p�vg`�s:��]���p�E��:��
w`tKt�ۜ�7a�Q��hT��VP�(�! �yp�M� �y��<�=� �� �aް(�zco�݇�c�lޘ���P6\���������ER�)BE�{�T* R�=���P7b� ��ч{�z���׀�)�ý y �3�^�CMOmؼ���yHs��(�� (��+��D�%UJ(�����{�t C����R�-c� Su��@� z�Y�� �tU����nw�����������D�UQΒB�
�c� (,96p���zCC�=� 
6�tI=k�z�׈��Oc���S�4:�/u� ]�^�@��u
@H�D�x�z�<�g{�U��� H�w`��{�{�{��B^�@��y4� {�\��rhEJ��E��� �
����JQB!�Q^f�wwI���OO{ y ���ۀ7c��3�� �� ;��@=r��$TT����HQG`w�����eQ��u��m�==�w� `�w;�vz {� ��l]`Q*	T�Su�*�	q���T]k�-�= ;�:(݀t� �t*f@	�����=� �ݏ@7 �6��r���T�)@*�2 J�1zw��� $ mХ�X@���������
(                               � @ � %*��� ��C&�)�0�J�hLL	�`	�`@4��L?L��	Q��M �d24�   j~E$
U&�#�Ѧ�� 0��&U%6��4��  �� ��B  &�h�jx�L����L����jmG�����~��� ��'�,���������]}Uς�?DD1�7QŸ�>�ٙ�C���m��m�z��l��s����$����=��c��l��q���������]���?���Wۿ�<�w�v�o�������ۑ��܇�ةj�n��ffk�[r���t��㊮�s�3r�n�+m�;��f�!e��G���7m���V�96a���w���7Ѿ÷��>s���i��};�q��w��x�on����٫6�S6�l٫cf�6jf�m��f��f�6j3f���6Q��Xlՙ�V6�[5cl���L�51�Q��c1�ff�6jm���f�6jfd>�G�ru���?���������?93���zO�|O��ǎ�N�����_��}|gC�q���f��qn˿�"��������R�S(��V��U�7�u8r��lCȢX��5b���"�L���i�Y��t�+f:@�j��Ӕ���XI���X^3�qҼx�#Y�Wa�#�B��nҠ6T233X��P:��ý�M٫��C��e��Ų�P�A����Q��z3Y�)7������ء���em���i7z�7iɦ�ޔ���X��5��q����휗˱�d������m��E�V3.�2�;Q����3�:�
!�F���d�n��؆�dj��+��c>ߊh�E��B��R�EPe��0X*a4t:�R��,���
Z�v�:�ῄ 2�&�=z��j)1�̵��g՛����j�\z~Aȩ֜j�ܑ��/֋�,ej�;�E5s��j���2�ɵr�!V�-ے��b:Uhkj�;"�V��,�7h�u�k9�5��_:Uf��i4i���{2���B�:�Y[�Y :Նի�0���	f�pI�����U�����J�A��NZWAZ���	�5�0��3v�V�byOot�1��!�nV�AW�-zN�0�f�B��1�t1��ҟ�Ǉ
vk~gj��K�����WQ�I��P%�m��q�`m�F����œIb��	�x�6�
/C�pEn�"d�-�V�ȩ�ǉ@�Ɋ���hJ�^���x��6�m��Ő ��Y�<�6@��P���}��*���^���nK��6%���6,��40�(l�4۩a�Ū&�02����/(I�f1+a�Ә���t80�f+W]Ԍ��C&��R8i�XH00��.\e(Sb����6
T�je�C��l��yy{*ˢ����ج�\rB'i�Q�`^]1{s4òm�B�A�������laܔ,�&��`723v�2���؝l����v�ݹ�Xş ��eѴ����#��)Jؔ��҂�&����ҥn&#�Z�p��H�5U��
ѠǕ��m���X�A�Y���t���u��h��(�Mj��}���ww�f�b�w�2�b8�Z�e�����R��q�e^���TLR��RVU�f�oE7�k��]hJ��.Ы��f�a��nX{���@b�c/0��Z�kU�c����Ad
�t]�t�0�0[�%jTd-��yYf�H5�B�ذ��\R�5��V^�	�OYu��F���n�A�i2�3��8���Q�6uO.h9y*�Gi���;�2	5;Z�7+/i��I�^a3r�M��^T�G$�w�U��f�X0�X�Q��Zݬ� ���Ӻ3 /��q�ێo�Zj�[N��8��6�ƣF�6ڀ�nmH���ji���A��/3z65�̠0�Bw#!���v� j�Ȋ7Y�90�W�����V�;:�0dF���1�� ��͘ƛ��m��p��kTw`��g\���-�b�`�"�.�#��l5�.&kk,
o�C�6�`�$ vڰ��JnK�b�8(�`��H<q&e�Fp���a��V�݅�����	�՛��f4���5^h�4���N�P��7Dph�6�sJ�2�J
++
ʛI��/1,��Q���v�+E�f͕��*YE[yN�Kɴ���)��꫹��TPm�rjF;Nk����"U��B�6&��n��i��n(j[�����F�/@��uh��e��Ǧ��7�]=bi�ս�l���y',Д���[��V�&���B
��E#X+���1֛��5Y-:���Y�c錃�`�����cd�jq}�]�.r褕�L١eԲr&(f#eY�ko�
QXO�P^o�o�(�t���1|�T�y��2��b˭�9�Yy��sm�ּ�EM̳�Br�$r��2�VDE� ���SS��3Hf�*�����5e2�[-��f�!�Rk͖]J��ɖ�I�-�Dw�n�=�6-te��0�/%Øe�X���22���$��ˬ�b͋�X.D[om�n[N�ۭt�V�a�5�[R�;KA���:\�Z��gm	w�1�p���ǶN��-V�T���B��0�U^`��%pY��Y/U`�CTQ�W�5�*)yq�j	,_T�l�����hU��כ�d��*P
`��f�;.b",}�
��L{�ЏE��k>�s`J��J���K������kTe��j���@�DSh����(]�fvE�鏬=E�Qʗ\S4� �'3L6��v�x�Ѳ�̩
�]��Kr���fU�:B� H�R	��#\G�X�6�h9j�C�ek+T'2��(S�wp2剡��J��`u.0�㼶wH7��+N�p���5m@ҫj,jTF�unU�wPa9��:Ym�6Fo*�]����2��*���nE����or}������ݧ�%;�u�(]���(Э�@�j���v�����gX�6��I�X����3P�r��U�:e��۽�,�c/r�v-�1��im��-�x%�x�z�D6�Q���Vn�^ڌ�w��Pm�p;Y�� �yGR��Yn&\�D_�W��>�2��3 ���@3#z�=�`l�N�ȴj�mUͭ�N��5��tZY��7X�PK�3p�������]��E�ؖ���Gk+��YnY�f���!�����M�3Pq��Qɚ�,��ZZ.�V��U<�Gr�U�ϳ �M�����E�R�Rn;�z��ۭ̩}��խV9�B0$�ƭ����$����\�Ts.��n���VH�w��C!��B8�2��2T�hi�iѭyk��v�ܻpe��sD�^�1]��vC��2l{A6w{��Zޒ�R7������C��+C(�X��
2g"�Q�"ⲢR�:֙�4t�%�rr��M+�(�i�/#�]ݓU�A&�;U(�Z1A�G�U�K���݋e�d/H�fI��=� d��ջ�Z���Y6�QG.�F7~G5vU˽�L	�71�w���5��2��ZE0C6���J�����2:c��gp�e^��h�5f�Y-Q�[�4���cj�-nJ�s�e���fY{�᷄�_�]��Q�u��u%�̣@m�uEW�T+�Z��&����{,��JӦ+�k�v���c۠��k��	�%�_��72^nc���v�Y�'b�7�JPb���Q��f����d=4�P����`�Ey�=�ӷ�!�XFR�6�����Jt(�&%̓���i�I������zv�-��������W���cr�:JM���l�����EB5�V�r�"S�`%I<�	r&�&+�3=S����/+�K�{�����ۦ�5n�8f�Q`�!ö��L�u�bh7Y kL��RbE7����]���)��%�[� ���r�h��V�s�J�mM��kH��1^ϯD�W{� ;y�&�)�2��J�2ٙp���)�ug.�2�,�2klS�̵�����x�1�����p���i^2ټJ�� �+
��]̫�7LJ�*Q*��=��۽[9��k%�1��M+`�N�ʲSn��W%�Xr��j=�u�$zr�cF�X����0���ol�̃�6�ŕx�=��o2�����o�AiE��Rf��0�˂h�����"_�n��fmэ��W���H��kӹ�h���9�i�n����<�&��$HM��Tc�34�C�CnಣZ6�2��������1 8��z%�z�n�~@#�SU<5G)#pᓅ�DРb���XBE�73��*0���4-��/Mo��`��sj@� َf�Cf�,���{���Ya�n&1���SzgbU�[�*V+t��O�
,;�,e*3wq��;�P�P2��C�wTջo�+\�y����6F`pL���!�s����U5-]�u�2\���Зkd2�՝]m0.b%�H�[@D��M**�!���YE��Ŧ�4�ջ@�ɪC�	�h��x!�JU�ù&�t�=���D���WY[.��2~f���4-�r��fd4��j��n���:����ے�պȴ��?�"��RWdb�� 0pÕR2��	P�Q�[�^��2��ˬ�lK�#^@Y�V�˃.eX���kf�Vs�$ˣ
7fb7�a�M\U��A�{�#s4�EAjn*/��ed4!R+T�hEb�a�ZE��t�2i�i:�մN7��R��bZ�Y����9SJe��^`�.̬"B5H�h^��,���q�ɘ�m�f��q�AHV뛦#���J":���ݷ\�AX��I��=�J齨:2:�js!�na���6���ӴS9(�4P�",�D���Ɋ*��d�hɻ�(m�����Y���L�-2��.����ȪJ075Y���}@�$�X��"�U��T(�܊7�j{x7��HƔ)U��^҃7,�����*��D�]��
�e�q���IHDЕxQ���.�C`�oAY��h͂��b�D˔�%�-B�JK;hZv��wI�j�&-Im-X�B1�j�nEWl��	���a���iL�r��eH�0��d×J2����ּ��<��
��Y��(�*� +Q���@�E�/`�Ԭr��Ҁv1���U�M��[l�B��:*܂��N��V���`�����ptl�u"��[y�a)B(.7b��Xi�&������⽰)����ys�]1�f~I��G�.�H۩Vl��uz�F�/1y����ɥX�<�R	!%X�V2,�8��w37U�BSQ44�f���������.�iֲ)^���D\��'f��m���u�e��1�4��q
����jf��.��Y��1�9c]h���Ρn���@ڛZs/Fc�&td�n�!��z��ǔ�w�!�ne��n��7
��;�kMLN�E]�� ]��4P�n�r�jmѴ7Qz+#r�3�]�P�7���p���ߦZ6F�T��=��म]�n�ԳXp�t��K  4 �2�[��zq�{�k)y�qV���e�5K.��Pb�·�ѴZ.���j�D+�f���.�4�h�6NfA+( ��o5ؠ��-�d��w"�h֪w�R,��ݙ+3k ��/N����ɗ���͔e`WVJ)���FI�,�|OזVT��&-MH*��Sbݦ�YڑM��bV�@��P�V���l�cO#�vj��6P��.B�P_Y��B��8]���dx�n�hĕd��w�58k$
&�jg!��;vn�u�ߢ�`�4����e���VVe<`Y�׆C%ƛ��xl"�*��p,�j��(d�>k�FVD� 3	�3灹�h<�.��	5Z�p��d�t����=�H�O ��Ś���̅�m�,t�R��n�+GV t7�E�tt�5�1�8򑰣����3�.��e��;�"ʘi�k;6f�LN����]A���b	t��̚�:��5:�lŢ��l��xK�w�&��n-'�f����.�+��RoeKC�%V޳s]�n�:��gIU˫��-Y�]횏2�Z7S'I�e1c"Z&\�53x�e2eҰ���iQ�b+�ً�Fi͈Msv��p��;{���v&�x/5pթ�MV��[z�*��Y�<bF'�낔f�#�@L����˺9�@X��M���	d;�Vj̸�+�P{��1��a����v&RZ�e<�+M�E\Ê�-<��{B�wc��]٬Ka�/n`a�ˌS%l�� �.�vX���r,5�[y�ݼ�o(7z�֦�p]� W6�cp�m���u�fh���e�����Y��Å�4˖-\��,!��j�(Ĺ��*��*�(:�G��fFdw�Z�Ǚ�Y�塊�[NHbp��[uVC�w�n�`��-bĤ�P�р]F�Q�"D�4c*N�(�˅��1v2V9�9��.�2�ٴv 7L�����M=���z �5ԢfjS,*Ĳ����h�� ��&%V�e�GS̘��0S��-<�ıI2��Z�8�4|b0H�.����G\����������e�x�Sl���?K�����0����f�?G�D����s��o�w������W�3���q�˹���枕�:�N���'�?���!�c	4P��.�k��5�َ��r�e�ۯnz6���F�$st�e��*Cq�\����۶�nS�E�u..;pܖ.�8�\^�k�z��T�pert�v\�W���շ�ή���4c�%�(��"��l۷5��^'�}k��ۂmv+K4�1,�P�4�.��Q��9z�]�<k�y{85r-Eܽk/3�l�Ѧ���u��vͺ�f����w<U�Dr�+�t[�/�r�wc]sWa�`�8^��Ц3Qн[�[�y�=u�<�d�zwV�y�<j�y�*�,�梓]Du���-�e�[���(�B�w��۱v����v���ogU���v���Z����j��BaK=K���sYrRj��c@L2-������*�Y[J��-�2A���m�R�Z���{Z�ʸ�ɓ��ٗۇ��8�=��#�K�6�裒��nIe�ґ�g[jE���^]��#"#��풺�V#����[UmV�ZنY�20qns̘,�PQ>����$���l���2f�66�E��Gq�'u���Å�ؼ���.{+�|��9�P��n�9�����ʲ��;[[���wn��EςU�k3���`:d)i�D�"a��7��Hʻ��GM6��e,��9����� Ѳ�M�\tQYg�b���N���\N9D�*��r�]-�@���ķIS��%�*��a��IG].���d�������<�.�r�x� �g�Em��:ym���.9uli�}�s�v��%��j����g]h���H�#��
�[��@�2y�<�k\I<v�]<��j&4n�B�F�l��4nX��GrKZs�[���ts(׀�#f�G@��z�vd���MCCMaD�V��(YQ��m�n��֥�J��dϓsl���w����6�v��H�f�x�|~s�o��ݫ]��U/lI�dۨ�Mt�m��r�5�^۝��ax`"k�3�3Ek0�\��(j�R��ѡ\�"��u�۷l07X�)woln^�q�݃�3�ᗂg���Ҭ�F��L���t��s�xi���7��ѝ�ưY�Q�;����Gh" �I�n�d�;��;�'t�vY}q� ��u˷��]�u۸���>6[Ab���ѝ�w�3Ì���/iq�,z%�Ĳ�s�j�,Gm�LM��x��2Z������]��E�/3v�z�4�l�8b�������s<ݤ��j�<�
ru���Z|o9n��ў�^�On[a���wS�m��P5��l`r����vS�g+Z��"J��GG;�rbڛ�᭹І���˱ɸ�@��O���hy�wA�s�p��3Hz�����vFvtW~ڌ����9T��]��9w@K�yv�ݙX�M^/,�` &�<��{0=�9�펽21��#����SY؁d�)��h��]���m#��݅��
x<�0�JCi�\�V3�{a��7g"��C;���Lh+��]45P��ޑ{\�Z��׉;X��g%�đc�]���va�6Yk5,�l�Ͳ.�xh]�-��c�� ij5��� �����7^S��E\:�ď]�<��`f��8e-�˪:<���iH�2:�2�[-�f����[�=9��=������+V�#'�m�B>��ۘ[3"IY���)�Zf�2��<�\m�q���z��]C���ǜ{��ꣷ"O3��I�9�cC��;�+��̈e�7�J���*��k�c=��f�8�׶�n�@����'�p5����$��M�؜
r�3��Ci`�Q��*T�eh���qȣ��qZ���.z��&�ƥ���E�7�-h��M71�3i�C�n�� ϸ�l�[�.ӣ-�f^1��kMl��gsvrs70�{p+]�p���ݍ�lI������5���6��f4fE�2�XMk\����c�eSHm�뒹��؏]�<��ԑ��lvlZ�z{sΘܽf�.����g�c�3�Sy�*����9Tc-a�i��u��n��C�m8����gM�Nv�����g��NZ-���a�Za����.@��6ۄ���]5|<M۶���F���nd�K�w=���<���dp%�5vw5���Cq�q�cX��,����\�.ʹ�ڱʚ��z���:|��V�L��n��;�ݷ]&�����g��^�x۪n0�p��๕؄��Ì��b��eH\tiE�A�8z�q�#ɎF6�Ǔ]�c������3a�l���v��7:�[�ܺ׍(�Ǜ�=os�gKlq�Ǯ8���X.����qk��!��[%��G��x�M�4���!�W޷l9��N��#�n��Wc��š%'a���QX��f�G2���ˆ�;{6�WT�R��h�s���;�vv�R^�C�w@���N�[��M��������3[x��t�Z,/��c&�t�
p�'lK4��=��f��`7:�ݝ㾵ɫܕj\dٖ�c�XJ�q����n+����� �N.^nǅ1�`����������y��%��`�Ƹ�������7c��xۖpV3`e�D��cu5��nӶ5/u
F-�d��A�UqC\�f{n��b���|��m��̖��U�.9a��zB;+m�/$���v..n-�t8vL8��^ݒt&���]ag���:�6ٙ]V4Є�1��J4�v�#��L�F�v�Mk�A�(j�-Λ-���%�mb���V��^���k�ۜN�5;�u��*2MF糏%îz�Z����ɠ 4ݢ��F��D������vN���QX�����fg��-WC9��X�i!���.���+�ۓ�`�5ۻK�/�{�����e��l����uKvm���Q[�/3�'T��7/�m��n�{w2v��oROn&㴨kK��;=z�m�𚱋�؜��=�ꥤQ�^�8�9��n�>7g��Y��r�Lp�Nv��y��ʢB���2�h��G&�����V��[Ξ�[�����[e.nh�r�F{\����2��\���S�k+@	��K��\�+e�e.��1�5�"�W�z7^p ���Qz�3V=Vkƛz����I�ѻݞ5���v���>�z��OZ�u�/��6�U�[�ҝ��/��4a�YXٛ��+,ŮՎm�y�<�0�r�t�<p	tF�-�����lh77���N��Ս�[���g�N��4QFf퐪ݸwH���L�m��p�$؍[t�����%$�>����c��^����I>me7	��桲�Q;e�wdS����m�|���9�f�n+��`��hF��c�GFdVPۗZ�ز�|l�#���S;���f"�m=֗���On����v���,�`��7,�ݷ�.	e�*3�DGR��b����c-��)��-��<зLh�ps�]d�Mn�M�ݚT��!mr�L通9�ݒ9�ݷg�<WDݨx��{��I�Mv�s���u���*0 ��и�4o3	���l�r.���L�ZV��È@�F�a �(M����uN�r�1��u�I3��#s�Ȑ�Zb�ɰ[��^\[l�R�ث��ZϫY�3�Kڸ�ǋN�{P�U��7:p3�=�2�=����2��JX<��nmk���j�ۉ�����ܩ��jc荢N::ے�u;G��I1�6VK���Sj����%�%]����Ga4�3b�=o,�fk��j0yZ�v����ki�)�77$�m��\��k�70�]�iqc=N8䎸�07+�륷*��\���be۷���T��8ގ�ڮ����q��yvv���Ɲ�;f��雎��qL�Ў&��cj�8�ѐ���Ѥ����ӳ+]�JMq<�T8��^l9��9���9�њ�+�a�)2M�\[t%���E��dRV�U�7D�87`��]S�t���#TV�C-��N�݉�r�v�pb�t���+tN<�^݋��ɺ!5�e-�&�5U-DK5\���]F(�戗 �r�K��p�;=ہ��9{l�;^�K��oV7\��ni��wj�z�<Վ�;h��Y�ۊ��K�d���k����v��7��nt�+�ŋ.�V���հ[��q�c�OH/O��s���y֎b�K��w����M�b�5�kb�X��g�ͻޫ�F���б����m�;q���=���iGGeI�/���uP5tqn�!�'\qd�D����+�8�mٳ�,ю�\�� ֦Nʓ�H�a+E͵���N�XJF��5���p�����O/Gnj[	����Jzv�y�Q�r�;	75�G6�����G�������1��A����#q�������f33v���O��y�v�v����6}����>Mo��t��?߯z�4��yy�
������,�N���yiU��D��2��lQ���u�|/�l��6�Չgs�=��Q[��Pg�X�	0$j�6dNኍ��Y���zb��Ou�W�8�3�<�����J8j���1XyBow�����-K���F�1���]3X�G[�8/+��J,�Jّ�o�y�K"�|����W��Hy ��+����˾�e]4���;i�� T�kJR�#�|(L��[��AZ5#;H=��)V�����	"��C�k8�uk޾�m�|d�`���W�:�V���k�U:�0����`Wf�-����.(��3v6>�[��)n��*C;�ݳ�_`�.`5�\� \3u!�ܱr�{��u�i�͋���.\:�p�xJU��V���zWv��W���ޡ�F�7l!���g���x5��W��v����_�a��J��4I �A��
�h�Q,Q������yN�<Bm�Y&�;�p�.kuŪ9{E�v�"Ӟ��e��K_K��T�3��������\�+������\�����ͦu��t�V��;z\�Z]\�w�)���uon5�kqA�7k�$n��m����r�C���"�����m�Ժ�+�`��<�oA�
*Jĥ�̆(�p*�M�i��n��[�l�|q�ǜ�G���(�#ε\��=XY��	ĝ�*��0)᢯A�E�������
��m���4�e�K4�c�l��	���ku�����V���(W�r�u�l�����+ܳ��S��m���{ř�X��>156Xs�r�v��4Uj���f��Gd�]�eie]0N�Ƞ�+�-H �P���J��=DiNp�Oa3pvio�s�~�R��啼m:#uN���]f�7��uB����Ln>��u�i|,�]�c���E���V@���zd��RTo����5�	]��yy@�,�z6;��[�cII!���VQz��h���/b˪�8i^��1\�_gp\�u�!h)�wl��Ӳj:\�f�r�:�]����v�l�^�Q��ocv%���5����=��X�N��S�١�,ᴬ��j��4��á�n
쭉�.M���WeS��wRK9�V��Bǀ�兠���[KXN|�urhdk�d�`�]�=;pu�Q�Vݚ�C6�-�ܒP�RDb��&^�'i���oQ���@�#�֬���+e]�t��,k�s��g3�L&���lVd��q�G���(�l�ch��h#,t7JE��>�JMB�b�0���s3mlofK�>�M�l��z�j�l�z��7�,?WRY�$*�>+)�ji��)�V����3��D�Kν�Q�ԥF�!U�f�r𕵄
�	�m����O��கk�YF���j/�;u�t�n�TW2Vt<L���W[��+t�̮��b�v��s%;�1��'
��H�B�pJ�菍mOe�u4��t��w~�+o�Y�,kAb}��\6 &�H���e�1�G/.�wJg[7M���]�i���¶�M��j���S9���#[
0n���aU���+!�C�xp�MKA�MY�G�Uhb�8P����P�VJ�Y�b]��|)A��̅(��%�����)1J�,Bf�j#�7�M��"��E���yT�G>�{Y-���m�F^��;�鬙��f�.�S���y���ٖR�@%����x�{Yg����PW�ʷ�p�sKY��{MvL����s@���Ȱ�oۚ~U8qP,8�)�dt�6k�-1��{C���;��^ޞ��1;o�(P3t��U`T�-�n7ܮ�M���ʜ5���*�f��lJ;P�l��$��[�4s0��[6���y�n��F��'+�����D�璤��x\�G1���g]�v�7Xl,�.m���$�}R���ϒ���ܨ�zk�Md�p�Ii1�����8;���x��a=���C�uyi�5���6r��<��m��j*���d�Hg*h˃�3"�P[Y.�#zY�G;`�Ӫ��x����	�h[+{���GP�<�3X;±nЧ�P���'�(�$A�Ӈ[�NM��$3�A�9�O3lc�b�S��5��a;�G���gmѾ@M�^�Xi��׽WdI��z���oZWp�����`QjP{�fK#��� ���Y�2E�L+p+R�;-��F���%;k�)RsU�so{�Y�k��t��\�|�;����k{P�p,w���V+�9�����>$�eX��76�'n�m��wB9���"�e,��U�^�nյn���5�Y��9�Kص�4upܾ�pS[֗h�L?>�h�d,J{2v�m��n���6vU���V�S�!���Ե۵oi�t�����9ܥ�����:J��Npd8ވS��;4���p1���L�Y/5�Jm�xՌ�eE��.��<�K�w�rܸr��� v�B�%&�NEen�?&�d1�=�5f����o� osti_0	�$t�]Bլ�;&_L�(NX1q�>�yz�ɦ�hߣo�R�� t��u���YW��F�L��{��2aZ��P�s&3��W��S��%X��t�����69V�ռo����jf�]]�J:���P��6Y�̚kd8{)������ݕ]�%*t
N��Qpݼޔ����G+nн͎�=)v�_R/��~����Vփ��n��;�\�b�|���y ]��*׵gfȭZj��lwJ��W�m�Ӆι���"!b�9���ۦ��ԩ6�0V
z¡b�A�s9��]��.�%�U9N��:��f��OUÏI��%f�;j��Ϋ�rNF�f��p֛ϖTVn���i�fՅ�[*N�m�S� &M���������L�}��,r=�o�빙�v;n�α;��������uĺ��5�f���D�7��h����o��`��ԧu�|��g�����VX��͉e,ՙ�����`E��V����Ԇ�U�T.�꩸�Εs˛�?NFdu�*E/bu��i�9F��%tj��ʩ���6d��Pը�T�-,�T�R'2`�qt�I��Q�o�}�2��|jont\��)��j�>�;��,]�=H�&�뀬���+8R�o��x�J��9A�)��Y�ٻ5���][7���n���l�vS��	\���-�h5mY�DR��.G�x70.�����(����{;���[[ϔ�:TT���faܩ�9`�Efl-�������;�&�X�jz�f�����,9^s���cp��OuJ^�l��8��r���:�m+�f��^����DQ�#��W��o�S5��PԖ�3r�y{����/z
ٓ�kM+��ؾT>�h� -���Dľ�/�^������9���-���N��|��-���v��DKh�C�e$��<�������]r;p�w'-�n�pY;�RLx"S����OXkyK����t����t;�������H�Z��َR����ݬ*q�y�>DKݾ��s�5PJ{��Jae�RΦ1�h�&ֈ�:�>�}��`�}K�b�֜���j�s��N:����W����� S��ջ�@&�D����
<-�Bwv�ӭ9v�V�ս�N�qKr�]m���:t���f��,)h���ݎ���|���A��H���[nP�͖���PFd5`gK�ۊH�:]���\\Ƞ	/����i]˶���.�0�4(���������ugr�쎭���N�z�J��m��՘�z�Yv'eu�6�"tP+��P��lϡ���Ȧ�2+uU-���J�ۥ6� ���7�nk��j�@,�~z��l,A%4����j��ʔ����E-
̕�uk��ω�Zmڄ6�0�����H6���`2/XӐi:vv2hV��1Y�n!1�O�Ci|�;ک�4pH�u
��i�wl���u3.�qV^��m�9Ev��έbH�5�*����I]/����ϕ�����Ft�rn����R����7�N���6�]Yk�`��;XoVK(�P����#v�bar}��w�E�f�����m�[}ۻ�����j�Y�؈��.ON�m��xU�x�k�[8e�'��]\��"��4*� �XjX�fǪ�6e�@�N�NV9;���;:7Nwe0�%ם�06ss�G�i��3hCټ�o�����J�Nst��h�Xi�x:�����5��z^Ҽ=4��˃��Z3�� �99�n٢������k1�����F���ھ=�=3��=8J|���!(�P��gʁ��Bu�͋�0f�WC�,s�$gW��q�VχK;k]�9VR�-U���`���z;+q��:�u4�J3%�`���`�VnEl#Ujm٨H �Ixk���U9�f�z�)�T@��H��w`��u J�[5��P����}�^�i47Ma����*ڕ`�a{}N�M�<>�ӥ_T��c*�ejTu[�/�qI�Ԣ�zj/���َ�!b�CM���&CLS�4��p�֖�ս�� �w��<��Zw�����;���H%�th�f�՗2Jh���V%E���P�l�Ě���&.�܊7��,Lg�����s���Vu�F=�A�Qa�b��b ���oR.^�F�����r�� �L��ņ�ݝ�ۺ�\�V^� n�ا����Eu[�&�L�6���V]m�n�PFk��2�f�a��l�I�؛�������]�,�bp5˺�:��Z��=��%l7�����Ry2gq.��fj�D��EQ&|*sK�r����,������ Ӽ��Z$�q�5��Z1a�)���>wN)7�d̪+C�s5��E����юI-İg��{���9[�Z�H���&�����ZV2��.v3`�=�e*MK�CFn�F�W=�b�2�Հx>t�f�����V�V�&h��Ǯ��Lֺ�U�մ�u%���e�����������B�n���n&${{g6��3�d9�\ዸ�n��l�R>K(������{�m�����xݼ��[�v��c%�b֌#+��:.m�SO|%f�t����h�K�a̰u嚛wt��7Fھ�����\QK�ø����x^�ur��-����zuh��zH�ˍ"anv� &J�c1\��Xؖz�wv�������=����1WF�X��fK���z���J�_�K%�c��n��x]�~�Z��vᜍmf�2R�DV`�J �\�Y1�E��a���*jy��[܏mpr�OY��YET�^�d���1T�yJ�8r���@��$�=tNF�M�-,e�Xc+N᝭�OG ��ZF�=xNɮ�Z��v��F�/zY����z�&e[REf�	�xE�{,Z��i�ス��������db���9

JŒ�z�q�%��*)w��'X�A�2]gP��'f���=�ց�յ|%� �j�v���Y��L���%Q��N��P��d9j�K+l;���v�-�0�i�+��Џj^+�7 �{6��*.�i��E>�q������'���7�����d��,5��L��4u�n�0�/n�^�8�ބ�TqYm��ERt�rD�en�emҝ8;�j��Vֈ������������/o.a��KT�M�7-'�'T/P�{��H9l��wTJ2J�
�;��������	Kv�HAwVNZ[� 엍�7[+��s���5
4��Mh�J�݄y���!f<�ַA�|��Ȑ\9�M�%fsǩ3s��1*X�!��N�ݥe��W�!���١;t.Օg�t�6qL�E���wg1s5��RZ������k.��2����:�����]xM��ϰ�޲9mŃo��.]�D/)�M��4&r\e�]
���s���Dљc�J�d�S���`��K�k*�V�MU�����%��AȘ���1��h!2'KIZ���J��aɧ8oB�0�-��(��\!^��7G$@a�#l�E�e���;���G�~ǭ�ݳ33Y�5���9>O�u<�3<��巡�v��o]���o����˟W�W��+�k��i#D!ig,v��Qwm�]�8rMָD.ܵ��uOF�v�˻�/<*�!���7Gc�rd�rN�eK�zw=c�����u̻>x�PB��&����3����b7+�C]Ab�fh�oⰏ�t�K���:���5�W���8N� �^��è1��\�[[f^En�lrgc�V��e��p��l�NS8:�v���x���z9��v���Pɮj�눽Xу�����: :8*j6�\�X�D�g���vN�v�z��m�H���ɝ��m>p���7�\����ˬ�Y�^F��|���f�k�1$����uִ�<[�B]bq����oWO'F�f�%�s{v67M���v�դ��I�n"�ڗ^75��]�m�����B�C�m��xU��a�z�.y6��g�	ݚ�nESe}\,g\�`���I�K f덫v�����"�.s�{(<��f�-����n��kD=��1�ȞɁ|[q[��wG����c��xg/-b�e6�'X��M������s�ܹ�M(����E�&q�a�E� jX�����e9f��Onms��U�j�m#�1�h��la,�ba�h�M�Yete��b��U�L.N]�M6]+ˡ/�[��D��2�e#s��+c6P�=i�f^s�s��4�kv죵�!���:3@�q���^w=t��@n�r��:N;_cA���8��f}zҝ�/*ǖl�F��!���`��[M�W� �Cq�l�t�w5��;q�Ѫ��G\.4�:�箽�����ogQ����k�g[�t<�#J�z��2mZ��|�i���-���+A�q4X���6�f�[��t/[U��K�ve�Z��"�/	tH�	�wy���`+�N[69��pX&9���r�e��݊5��R:Y"9-� u�Z`t�8�SF�p���Ȑ{j���D+#W������m��}N�R�ȹdV�ue��*{xz`wvSPq�;]	.2K/u��$Rn@yl�{�a]3��̉,*��T���()�F�q�L�³�i�U��&<«a�7;�a�+K#����j��"�*��LZW��;��xm���d|p`q�2�VC2�)un�	�����BT�FcV��l�Cp<�5\]�̬r�
�{X�9d�mq�0�$��<��5��{�{��i(�-^+8E�$J�`�W��{�u�qB4wCQ2%H��ع:L�4�hE��
I��`)4�(�Y�	�ߕ��@&rX�CM���[X�������I$�1��]n1�c��JH�S1���t��V��C�t��̡�NJ�|gM�6��ո� ��H��ѳ��|l��Oҁ;i�X밋��uu�eH����6�4kL8���{���f�JW��qe���%Ҵ��ݻ#�U��چMk�����{��9��9L�˨�b�2i��v�[&|F��kݥ��Jk4��)
C/),��@"Ƴ8�,�s])�U� �,�H��׈D�����-���T���p������k�F���v:vph����we	��nW�Wj���5���a��pv�5�Z�k��{��u֑k��K��G����!<���i{Kt�~"l��ّ"����֬��o_�u���X�Ed�U�-�l�!d�TA�8�U�6���������$bm����,~��2�h��<�S��S2��f��CV00������e��_o+����)�]D�8�M#|��� ����bo"�0Z ��*��o9�U+���@��+����̧�5U��3k�h2�P�d�-��I�X�iU�E�+;Us�u�켥��,�px#�YIV��0��:��E}���U�����˴gf�1��z�=<������öZ��7r7!�h��/X�n�NV6��;[�vtu����[��1g|�.gj��y/M*C;Up�#�u� �(�!H2�p u�#��5��� �\M�H�a�t���]L&��.Ѻg3�z"_`q�J_MT.0�z�D��q.�Q���㒐a�Ne&,�0�>��C(|�ܢ+P�X�.��]:S�U8�*�q���I@��U�y��@�-���=�R��x,_AW�ל�*���i�`���ɸ@�a�L��Y�#8���d\I!�Q�ʬ9B����E��r$��1CY�w� �M�tW���E�Z>��찰���5ap/%9p��D���O��A͍�GiD���A���nn��D����';���&���[D��0�L�bOsRh�s�����t��P���]�N>�*9d�h�����h��p7NJ��s+񯪊X�}MA�0 2�L2P`\���#T�(+��gl�(�yTI�9)�T<�� �������PC&]
�r��u֖��2�{!��^�;����ҍ;�G.��8�n*6^Z:m<���;C�!D��yV]�F���a�L�~�!w�&�!o��A�L�I<"j(L�:z��og��#s����hsk��KwO[pW�`��L�E����2��}��f�♈V�LҦ�hH�!�1%n+ن8	��1�GF5m��l:�[Q�Cf����gQs���j;n�����ߟ}n���2�U�N�W1�� k_IU�)�&��j��2�!��*"W�sMQ��{ԧ�)ΚTi��'Ġ�.4�l&[L-}�����!?��J4F�qMB�.&Te���I����"� ݅-����v�{����,�x7�Jph�O�`���(�Y��7 �]i��}�v��G�R�׬v�}4������ve�o�Yx�{2��.G�vd��LP���JfD9��C1KrX�bx:����
b��V��C@r!F
*r�Q�'�l�	� ���ݕ/`3�LLͳ���QX�uTB�!��t���n��v��
�kyfYu�z-zt��۞h޳�$3�MX~��7�_����Jߋ����2�nN�����=8"�fE��@�o����H֘pSh�Qf�9���&��h�=A���0�z�1Kl
B�v�8ذ�'~��ٲ����L÷��� E�������UA�6��EC"m��G��t/��%3y&��.e�q�A�0��i� ����U��'�fG�h�AU-m���q����l��JDe���U��|�RU��� �{U��jfS �Z��ýJ:��ΛY��E�:�T�+����2l�
8��x��[k3�R��Uw�]���k��P�AК�|[G*q�7`��ۋ.��fZ���f�ds��A�+p���']�k�1��u��6���J�G<a�C�ܦ�۷HS�ۀl[d�7��,d����� ��\��q�wPgs�:�v^FZMj�����z;�|,<� P��?*@�B�m�����2˄����bE��	�m6��x�v�Y�^�ᲙѱAvm��ƚ��}3������m�~C_��rj�/8�b%n-�"���
 Q`c��J��t�(8B�`�n���3�6�:�S�ZF2�gS����0��껑 E
�r.�Ӱ� �N
��eI��{R�U�Gi]�'����eT򝲻&t�t�@���
��1��iħD�Qo3Tݠw��2h@��yj��ky���$�`�-ҷ�j��Dp�4��6�#����և2�/{\mW�$�`� ��e@m�暔׋�) ��]�3�h���������J.u�������z��Ǹ��i�^��+���	B��U��<e�e�a%�њ���Nv]ӂ�X�Y�FU"��	�؂��:BFI�@�����jQf+��5��,��(��t-�ux��jiހ���|�'W����1�C�t����(��C�Xoh�S+aDQ6���]=�b�\%�h�F�^�����i&i�����&�z⯎ԥ���75kT�w�(0�h�9�hL�����6�"��N̊yl�35��ҖGt�&9��6Z����.�����"��N���5�����;:�v������@��_0�[q��ڐ�r͋;W���l����u,M�JP���@�U�=f�6X�eU�q���"����2�b��LE�H��-��a�n�k�9Qb:��Pc#/^�#V�΍Y�C﨩o�nŸ-(i� ٤�>�1&ռZ���4�Q$Ef6�}0�"q�8S�A�Sf��w���pH��j�i9�ЫgZ�ś&�84�I�P8�X.oK��OR�T����0��*Z ��1�ާ((Rb��[y�1�S�j�41�}�����jg[{�
$ᔚ˴"�gY�p���qpĪ=������1�껳�B��-�UT���&�H�E�J���.k��<.�K3rV<�U��KzT�����=����=`�
탍�0*�K5]�g�l[7	���qy!�q\.	��Y	�&{���EgN�A���v4��]�H��%�x�8b�Ъ�EX��u+3n)�wP�a���om�<*b���񙂖���0��0�
��=DM!��Rme����U(Ż�z��.虁��p	o�HUp��KJz�U�q�-�U"��4G,�#����<�'���m�r�#(�
aIae��0"�ب�W�}�N�8�9FP��_v��(Y���D�(�,(�	� _q9V>���hڢ�Yo^p�wO&��Z�1�,?�P�qX�:�K3�z���EoJf(�{�3F�?����=�Ӥ_��z��i��X�5v���P�1NH����(*&�f�L�ᰃ �''L骊F�v�#o��J՘t7A�z7��$��f�,%�*Nb��f�(��;v�Uqɉ�Fg�UwR�9�2�1E�a\&�$s:�F�E�6r&�9G�Ҋ�_i3�S��!P)��&
a�ٸ?]n�u�������.��sI�v����F̮u/+#%A#��H��IY�]��nұn���c*�̚��5K1�"�ێu�bo��(�`Bޥ�@+����V�EG��&�暠=[tK�+%�M�r8��-�6�S�,�ee'�]�����šA2�'��f�2<��̒G:sp�u�n��jJQ�Ѷ�m3И���O���b8L�%����D�����&f�'���t񆧕�p]k%��#�&�6�8�#�Pldk�ŸE옟^,��{���7�Y���p�մ�
���nx��/0�q��n64��;�m�Tl�
�Q�.�(�H�φV����tv�	���,}c,��N�-C�p�I�#;�ŷ&mԺ�J�,�bKm�ŏ.��z�;S���f�����s��a#����y!q��IP��7g.30��Q�(&8M	tP�{C�RE��r�@޸q2PݝFֽ[
�c��P6T�pr-�	�	����1ϙr����7��c�"_�(�4,*��F80�i0I!!4���y�p�se��2P�Zq�:��+���U��y�te�e�0�i��/��Z��|ǟ�e`�����J�����=��϶w�Z2���m��s�س�\]9�E���7E�8���1}oEc��׬柮~��u5Uu��֣Oo)a���	t
5�����4�����9z'unQ�jd]�#���>�[e7=��rcj%~1���ѱ�������_[�#(�̲9S݉f�TЋ)��G�x	�W��BN�An��P�է9L1��V�>Wu�]1��7QP��y��H���gUE�U�٦��|�#��P�B��)Ҿ��wkk�|@�_E �j)@��2����@p�&Fn�|I���@\��j�ӬX�J3`A�&b��q��8���PT�((�����AY�;�}����ai�5B���5i�0�u�{`�i��v��x�1�Dڞ�����f@��h�j�oϾ���� �7�pIe��66�2N-�[v��6襠���9�� (p�E0&̣ѯx��D�^u���d�;��M�ә;F ��&��6���p�A����d��O+�8A�? H>�߷���7�;��dѨ'F�q�3wmP_#�E���:=L�u������������l՞�Uf����1��n�,�-��`|ǩ��Q��.cz�E��`ofK��E��-
ږ�T��)�^��<(�jp�V2�A������&��GE���N����n�8/ ȦQ�:��uh�9,N3�,*�pE���ۊ���9�]zT��#m��u^�!n:��i�!���3���5���6�'���Z��-�W	���j�aȩ�����޻>�u��mJub��y������M)t�rwn}�� >�S.-vf6hf�V�m!ݞ�E���ܽ3t�����r�Y�e���n�7rr���,���VM`7�L��d*��.w2��["�Di��0�g��lJ �}���wg%,���1��dh92&�`�Ŷ����TAv�v1��*���yO*w���������qԓ��P�-\�푔�n�� �{[��W+���)��c�ɡ D���.�@�^�x'��r���i�Y-��ly�/:[�S"C�6��pc[6;�ոX1ho
''vu���N�ǆ�$T�f��lC-�����zo\�����`٪Ĕ�f�*o,#vd� LKxN�]E�~9�ĕ��w�s.�Ϲ�Ѻ���6���:٣�+��x*��f]'�F��<&P��%���=���5p^�����EݛyhT���ֵ��o\�F�,�-_-Q�}�^5���_�"f�x�"vpC[������2Sњ���-���7H�i����'0]�:����}�Wqb��u�h�9����{�DD��byw��E^�+����f�Yq��=Ǖke�[�9ar��v6uV,�4��n6�(E*���d��i�!}Q�6�>�L�ؼJ.�R�^����͇X3/5X��s �nQ�p�P��F=s/#US9�i�b�DE	����n�L��[�����u��Zh�G	e�����X�yO�a͵������|	싓k�vƄ5���	Ax�o�Iâ�<]:������Ǧ�j���!�!Gtn���CIՄd���ETX�s�)%na#0�Ct�� h���BF��р�1����wtN[}+r_b�wt)s"�[�.ux��)=,�[�9c#_ì��w�9qIM@Q�,T� °d;PX��l��ܝz�ј'G���n������mk�X�%��Ա��2���~�����}I�J�4@�
��X�������������썓j���ƒYBP��w����H,#io�� ��Dg�#zᄃe4Ju ���b�M��ƞ��E���%,b���q�H�B�;s�4�ԩs!��ݬ4�`8�Zq=<�}��P�&;��qm4�q��}��-�W9RM`V]�x$S���_j�:1����n�e��D��H�G\�\W�i�z�q4��_�NDRV�6�'k�ņ�{�1(g���u��K��	�2KXe���tէ����ٽ��Ƹ��Nrd����қ��Ξ�SI���YH��-���7,c��]�?ncz,��z��)�[�"�:�������xrS�OS����vuó������=��/���}����!2�1<�.&1�6���4�j`-=��k8�p���:���R
`%�S��aH�J`CB���т1��������)#hbOs��1����|����w1�kM��@�S��;��-4�I�Sǭf���Ȝ����
c�l����ѭ�JD.�b}}�6�IH��w������&6��ګ���Idu�ض�N�+ܼ)d=�1ݒ�1����K��\�l���-�I:
c��x����ح��.{ў�"F!4s�����1�D�m�b���R�9��5�w�c�U;z�Z����!`���'�<�1�Y;�R�&nl�47mM��%�z���ʸ�F�6����g8������.�lϽ�#I���"��Չ�H��I�:��������+I�sb�K���:-��z�
Q0e����_w�纘X5�.�kQeM�wm��F�1hw=�d�cL[O;�\�e��{>h�����x�]�SK;K�yW�be�*���v�ULظYy9)���}����~�Y�;�B�b�`�}�U��b�`�[����!,G-��X��;�4�jw��S�����5�vv�i���Uwa�iL�g��Hi
E-����Ʒ2�G��br�PZ�,�mw_np	cl���P� �|u�80�u-���m�=i]�}�A��4�K�}���GX�-�w��f�)�4��!��}@m)�m&%�r�������Q�6:`�F|s���Nɚɸ�Gп_�x���n�ENc�%�BX�{�\q��%��~�+�b�O���~��P�,}��^zק�� �T�񟚢*��WdSc�^<e��;B�����G�<n�I=�-m{�U��輚�L�E4����� (NP9:�9�Z�X۵�ܘ {m��s�|E���7(�.���Jn���`�Y���h��.��C�G-����X������Ͳ�J6�1�m�=�ܫ��;���۴���s��N ��9ں5me�����tro]t;���u��m���\CRV9"���ZE���u����:���_>{��?T���+��D��a�!�-�N�K8��w[��\���B9V��J�U�b��R�t0�6��2WW]���[��Nz9�/�.fjfG�����&&�3%G�?�j�n���s��V1�s!{�}VoG{<���,,,AlA(hO��;���m��'�1$���߁��e݇�Lr�o�ʳN��R�u���lG*c��lo�ל��%��_g�f$^��B�{���6�3�=�h��
 K�i���vK6�wwXY��M�i"҆/�z�6�v���w]�4 [�X� dȫH-�`��ˎ1Ħ�����d�:bF�%-'|�{˹�V�nWyYw�#�\���+��4���f�V#����o.�Jb�l$�:�1�4�Sy�s������)�ߪ��:�S�c���n&��f۷����b�i`��ՆݡLJV�
��8�p��,�On���Ű��{��9�B�>`�;�ɲ"S)5l��|�uwL���TYyN��``�w�]�2�;kc]�e�ECZ��=��ִ��7s5�X�7L�Hi	clGެ,Ǭ�n���긧l�cﳷ��{���Du��d���<��s�f��Ķ8�}*{鹦�h��r���q-��C����8�������9��
�y1��^���;\��},��`<5������� ���YV�y�/��+E8Q�>��*Q������Q���%.�N�z��O3W�6������`�E�!|�U�0[(^�1��{�c�M!��"�}��c�r5ٟ�[H��)���7d�\��X�uq�i�z�����4ű�;�ܔ�U;��S1"�
�v�֦1���ޜ���"y!m!�~���ۑɭ�s���]'�ܞ0�'^�j4�cihN�9��l6�$S��6�A�I�,1��G�{���U#�#��"[%����m�ؔ��"X�wE�H�)��g�޷��� ��Si,��XrF'S�>�G$RncoR/���ɏ�Ys>}�Ǝ���8c���z�&� U�W�l���[��t ��C-�2:.�f��*����#�3=�ۤ�im!����4���ض=�e�v(�uf@`�4�1cz����b1���'�uV�SVhʫ���G)8��=V�̈́D������g�Hbm)(M���\i�`���ޫ�N�o{�A��$�iP%4��y�O�tԵW4Im��������{�hJH��j�b߾~y�<�OPm~M~뭡���qjs���r��O�!P �hC"+9�]F�&*���Q�+;a�ڦbG=�{�)r0/-'�j�q�s�)����J�ؔ�s3�&�g2�u�����1(��_;�d@��z�VGQ���}�u����횫�ګ��E1�D^�=ꏯ|�RDb��٧Lb�{��q�X:�Kb/��^u�11�ͷ����6�CIM1���di	x�dH�MeI>��*f�̺��i�����j�~�b�;b=��Ϋz7[61�8�d�>��Ȋv����gr��Ɍ���#���B�00��.�|����мa$�iBAAW����5�)�:�i�i���`�oـ������سF�i�ɸ���#�Ĵ+=�VRi��{����% �H;=������ns�9l�bc��~��'8��E��77R�7����1����������U�rX�XlsshO&5��l�$���R7���cm��s��7	&�߲��C>��;�C<�J\��Ӄyv��1�� z��ͻ�"[e���}:�'$�c
n�Yb8�q�ﾫ2�����뽳LC�lՌ�봢���o@�dٴۈz����[�J��#Oɦ��U��iI�� )��`�}�M�4����e��Nf���T��Z�V�^R�_�;1O:���L7V�1�p��N��Ffr�d�PP�wz;�t�G_��7Q_�./2Y�D�P���aUR>5�N�n�������+2���/w�ʳ��ʕӾ�+wqi���i#)��~{�KT73uq2�Y���ǐ��Lb�ʰ�%��-�I[�sACHy��^��cl�_U���LBť�ݫ��P�&9��C���N�v)+�-�Z�n��]�:�Y7kaa���6�iK�I�<�sÅ�������j�s33+ ���-%�s�J`�C��B؊�0_��o�O{���b!`:�د_*�)1)�v~���M�9L�Pm�%1ʉ�~�4�nز�6��&�!]�����lsךr!lmNz�di7��h���!��1�n?_����v�i�=�$-);�{Ց�iO>����ȷQܙ��0�{��8���6�o�a�"�4�I|��J��qVV�2��+��xQ�k���t��)Hi	AJOM�ՀJJi�v�����Rm�>���:b�$��M}&}����V&�ﾼ�iĎ2�W{��%UYm^�������>�/�m)���B�)-"^%1W�Ջ1�ɐ-����#I�)�����:\�J�->�����ښd�2�Ҽ "�Cӑ$�jԒ�� �z�ƘcA�!;����ί�T�J.���A�R��ʁy�S>e�XFv]�iE]�z.%�6ӂ��6������f��1u�e"ٽc�9� <��J�3�Ky@�k��1!y\��p֋�3xzI�1ɪ67V��.N6�m^��6s歶F'\�]Û��׋��\��&�g��)����m�!Aч1�6��W�Z�#����7r�[<�˦�Mw�{��)�b^h�9m\&�J��
��T�TJ_��Uc�j� �J FR�0�8��*�ʈh�Z^M���N�AJ��	4�%�V�!ɸ��:��C\�^k��y��D�&8O^Gz���ssuu��)��	�S��M�je�I�e����G6�-�z�Ѣ�/��Pi8���B��X�����il�����e�-���7k��LNR~??|���/	��#��"�P�{5YO������S�;\�Θ�lc�����%�`�-��K�G��g���W�j�/#��9���3��X`Ť��-����JJ�&awxF�Ķ�*}ڳP�Q1���l6�`��Lc>�N������f�' ؖ������k��h{����~�o�H�!��e����w!~�ݼ4�H8���̝�ʮ����ߴ|��;|�1>�$�-"-�P|��İ|��~�4Ű�2�{#N��ֽ7n`�6�З����jci,Z}���AJcH'��7��s��h�/-�����sa.
�7�e�j��8������K+l�[��f�ʚ��&�@�g}��'`�[��Y�B���y�X;�w���B%8��
��C8���{�r칖�Y�eշKCl�����=U�١���Cӳ��iדKEh��ø\H�sY��`���ß����go�OM��^�3W=[ϩ�ÍX�[�q1=ݡ	��F�y�}t~xJ���l|b&�����g5���ƍ\��ƻw9���B�)�R����JC�}�ɸ���-/����N':Y�b�a����Ci����ns��m���"z$�I�����,Clv�����5��沦#�	Ԟ��m��-����61ɴ-���I�+u4V�o,6ı����7�����[������hRq��o}�o#��%^%�~�U��lJk�]l��U )m��M��؄���	��f�+2��4�1��\i��������ڭ�����N细`��ls����iLm#��͘�$i-$۷2�8�����p.+��ֶ"�&;7m:�510�!�)���$Su7��j�fvZ�3�fe�m���1~�ՑI�i�wrv��Hm%5	����q���߹z$,E1��$m=�l��������{Ws5ut^M�a�Ri���w�Ն��WI��#��B�S�v��LS�܏���Z;�>@�1���G��-��a�[�1�W����n�.�'���C�Ls���֋4�t���9��m�U���Uu���%)*1�>�rR��PVV��0D|j����[�3��xTIUW�e��T]��zwbx��i����ҧ�5�]<)�
�L4��j&j������Ҕ�U�ٯ�W�S�+��ii�l�1��4a�
Cm%��Hm�clE}�/��7w%T�sf�lZHo�̃HJo�Ƿ�x����O_�X�b�|�����i$���u@�;7cz��J�|ϊ�YE�٩���G��}�0<1I?r���wbRk۰�%8�BP�w&�1Z���~��'S�Y������}�~��hiz�XƠ6�q'em�FA��*�<7e�;JJ��>�&Z�z���[�*V�AԴ��ĘN뺰�lS��`��j�]�F��#Z$��̔����Z
Gݘ
`)8��3FDn��̗Ҏ�����Tծ�n�8��8LG��6i��{Sp�m4���g7�ޣ��$��Ȟ��ك��-��}�lci0q�p�#�ʁb��'�<�����v�]<'�x���3����i)����dD��K�֘%�%�Mz��bKClGo뛌B�46��4�(E6~*�Ne��0}�f��<6��)M}�U�!�b��'�׬0|�S8#�>��X���po�?g-~[��6G^k�[�=��hd��r�@�?Y�Bv���2v��7VA�{=��e�T��]�ȣ�E��l#�Q�ٙ?E@�-��&�8�H�j�p^@�i`x2��F(I��ш�4a����	'�)�~��F���G�m�ggx~"ӿ{VbX��V$�7���`�)��ٌS[��{�u���4����$���'Io9��?voٴι���vn�<+8|\�s̽�a8	����D����o�L�ӗ9v`�8�S�՘�'FO����bKc��læ����I�f��S�Rk��1,i�'\�3�m�����]f6m6�C���p��[�w�%;���`�|�:��>l�Ɔ-z�di)�m"��U�$���w�������'�����c�4���w���\�����04���ش�}�IM��^�|�İ]�����Nw;��M�b���=���hf�lf�A�mm��5�׈� ��{ �E1�l�v���L[���$����q��o��ޓ�s�~��F��6�^wU������:O��K%��yvb��G��7P�1,uf;����y�HJAg���0bS����g�F�w1�	!	����������w��V�z�r�: �Mbr�*ܓ��c՘b,(�x��O�"Z�e��U��5,��W�g�w��eq���%�B#B"���E@�ﺂ	ǩ`���FW�:ܗ�034(�����E^�����ul�A�
��� F�F8��������L4�]Î[N��q%��_��T�V�GM^�kWf\J����dgmi�P�񔴣��X��(����m]�mx�_}����6b�v�k��^t��f�y\�U�s�&N�0�����/O�u����j=&\ ��y*G�4m�'7f�9v��l�K�.u�z���i�ב�x�c���v-_�P�f�n��5}zF���XUgW	���xL>���
�D��u�8��_v��2�`ƭ
WY��^�q���HmOqu�O(g"���*�[�b�'�{Vܯt���+������xs.ߓtq���N֗��c�~��喬Ԛ�����85��s6����V�*8�݋\��0Ed�7sook:�onA����ν7Jܕ����\r]h��]�Wu���:� ��ڰ��ϳ;��\��2�:��g+���\岷wU���!��<G-݇��#j۔�Ĭж�~x�	�rDѹ�\�g]�H�TH��GP�;��/6i��+��]��x۳3��|'L�N�t�A���)b�[W������S
	��8L��t�9�;'�:N�S���m�to\mUy�G�T=d�y��J��4����<��7-����#2�4��˱�d�l*�Cxm�:-����E���8݈e��]鬠�"k6�X��2��5��������ܷ���k^
�a|Wxvi޽�g����ġ[ݹ���K��"�\غ����v�;r�$.͡��x��U.��0X��܄+l�&.��Cdc�ݮ�Y��ڽ�v]�
5�a�{^՛��68�ƅ�f�=�׷5nr�+G=JW��S�P˷c���o�a�6f
5厮�F�E�Ѣ�u�[�:�򥸪J�ʩ���ˇK��R��-�9��z�=t5>����$Fx�9��w�7^KRH-�
wc��3��L��D�l	�Ɩ:�F]Q;=�F�;��\bT3���Z_n�ׄ�z��neB��ʃY,�벍Ԇ��5��0ca%gv��{����t� M��3ܗ;+��#��<�v�vݹ尞�ë�r�j�v�c'o%�ѩ�b\�@5̪ˤ1�)2,6U�L�W[e�����F�����r{Kc�޽�L����PM��,�]��%�9�d$�>8���;���o>tz�nm���j�sKHs4t�n\i�UUW%������y{v���1�͌[ay2Mɺ\n��m���'�Kes�����+U�8�l#M,��]�lY,]Fk�2b.Җ�a�J��E���B)�H\���w\�lM��,u.��ƌ�W I���u��/\:z�q��n�kq79��"��W�ۋ��ƛ�Ó,���ll/2`��ns��QV��fV9'l9�*��&���EN{]P1.��m�h2�1�N5��n�'Q1����i����~_���2��s@�qXX��{�M���$\��{�@�����W���0T9R�z�u�).��?N;�glޜ���n`Z]32�fP��w*�&6d�r�N�,���۪�^)N���a�yn̨@����]�߶N�����T��DԤn�$�4lK�1�Y�j�ɺ+o���	E'�h��z �@�7��@��PۈUnc��x�ou�:,I�:7F�������q�4b/53OvpC���u���0�dVɏ�P�쭝�j���_��j��r�Q�q��@%P�b��P���!�7'
1n�u�.23]�vޖj�)N�:6I��s�=a�1�5�����|�T^p�R����^nH��C�;���Z�Y�LO�zT�>�����[R��Ng����Wh����e�+��J�z-��X�V�oU�g�q9(}�f0Vo[��+V�9weq��\2��>	���S�Ce�M�4�0��\Y5�HPgJІ$���Pa�˰vCS,^�	��w7!�9�� ���� 	*��A��9��*%��a�;$H0�C��\u���u���Z�u���*�9/Uf�ݶ�]�J
��=����x<s�Lm���t�u�>;onBj����tx8�7�8מ9;[�x'F�n��e�xs��T
��M*�ۥ��K�l�0<�B�ۍ8���A۶�Q�B�b78vIt�A]�ۊ�x�T�Vvj��3u;�M-TL
�\֘�@�l2���b`�R�p�{/��7wSѼ�l
���U9�p�s+/K��<#��'�A��G���1R����0�~-9�u�ӹ������w�͚Ф[��3�ꣿ���0,���'�N����LG�[�6��Ro���&
)�X'.~�p>�'� ����w�L���c���-3�I�1�o�Jc[������LH�I�g�"�-��|�'k�D1>S�m-���l��U�9�1i-%���l6�KciH�}�d�i�{���o��{��[XPRjC���y�6�LOo�Ή�JK`����W���b#�}�9j7Ӛ��
�Vi�H�5��q��%?'��w8m"�Sz|����|S93
)��Y������(�}�D�jn���Cy��B�6�i#|�yb8��/TA-�{׶�%ؚb�������p�bP�wE�6��6�$�O�^�r���� כ]vz�q��3�9KWVU��7���k�l���ಪar�tKd�V7xY�l��9D�1���p�M1N����Guʍ%'QO��6oA�2���VLL�䕯{ׁ�I�y}����7Z��I��I��C���X% A��'�Q�a�4va�c4���y0��|\r_VTL!�����r
|�u�W���N�S?)��z�DN�����چ͋B:iJ:ԭ�r�Wh����(��oVb�(Z��սc�1"�`�5��M�(m%-����q`�6�;�Q�"��QT�ۤ���۩��f�W��8��v�����z���`��}�<o�j�O�i�3��Y��6����s�i6���,�a�S>�������4m�B���Of�������y��#io����u��R�T�c*O�ڰ�[��]Wu����H'��	�&g(b�����ۻ��[�j�/#�JC�מl�H��j-ƫZ%4ı��d}���Ф�g͙S�2�Ns^n�!��Cl��v����	�;���Wb�ֺ�B�kVڶv�fn���`ə�q�����s���MP^�,lƮ��	I����l4��%��w>���)�E̜��[ϽU�%��`�I�1~ު�I)�-7��y��詹o.���,m��,ǻ��~9�b�<@���_7��i`�l_{��]�oS��\Mw����>�	cn0;��Q'�Q����Ѵ�lE�w����H�[I��M�N����W+��T�3��D�P	�!������VH��
$�ł�j7U�_n�"z��V���0wv�F��X.������_C$���}ua�e��Dԡ�D�PBԤ�%�?d����;^�x&�U�"ү~��sT6X�T֣*���ORS�i!JN�^����m~��;Lc}����l��1"H�j`�?�lLｼ�iv�����i�j����p�cII)�O�i#Hkڜ��ˮ8(q�����1��.d�=����6�����y�"�iIi��>��	I���N�ٲj�1����=��l�%����15�����϶����z��˹.dfkI<�C�E9��Y�LbH��;ϻ��q#�L���}��+0��N0:����Mvs�m8Ŵ�`�f�z�|L�SN
f���#�"�o��c���;��M&�B��}yI�)9�e��^������4ƈ���s����
`���h�յwUv�H�Y��#iLO/��_�������N�҃���q#�,���l��@�ln���/��ilW�wS=*�鹪�fVa�i)�����6�eaaB��Xi)�'ȉ̾�Ƙ���oOdO�".� �9Q<�ދ'**��i%��R�^s�?��� ��bZ�\�D�}!k"L��E��A;P0�\�}P��==L��>:��XH����B��:c#mKZLd�d:�B-�V1ʐ`)����-1���O3�s�f�J/.��8�8�BO���:M$�[<��q�=��$��������R�wW��+�ILN�wf&�z���2K�sI�og�,ZK��҆��)v��k"��;�ڞx:z�l�a��;" ��n�j`�)Y�ˋb�)9�}��;Ha�[���[.�����w���r���4 bB�n�-)�w{oHiӷϘ�jg�77����m��-)/��� �^��#I�Lm��pm-�H��l�/�!m9߻� �p���q���NT���B�[e8痈p�H��%!1�c�C��??��l�B�{]�a�-tu]�栎Y1���f!�%6Ŵ�����-��X�HW���vU�e�:˻��S�F��>�՚B�z�1���u���io���7N:I��w��BK+��R�j�0m�����$��̒[3U5f��i�=�����!9%��a5t¹1�Rw��[<�8�\���dm-�I`�_�q�-"�q���yy�ۓW6�m��<��A�����5G ��L��Qbة1Y�q���2����W�oJ�o2`ɘ�}y{T�4�M J[��˂.cK�ƞڵex�-�7�5�ˣ�j�D��]Y&3<�u�q�F_9N6C��يi�5���洙+3�r�2�;�cG�㫈���n�]�\C����.W$!�U���C�\8�x�t�x��,,\kwZ�=U*Xy�n��c�R��<`��LH��(��ʔu���Y��7�|s�s�516♒X���"�J%�ѫ������fP�,�
��4�ط�`�B���
 �D����A�ڌ�n�0H�Ҥ5�<�盄ϓ�EH�ݱ�xs���;W�������s�7��6�>���Q��Y���\bP4�_57�6Ĥm-��2�剶�ʫ�2�;V-'�a�|<K�%!�	b��"����1lEnA����H�]LW�����ܱc��s�a���KI�}�ƚ������T��BX���ٌbv��s�\Dُ�{3K����]�����C鹭N|�S1�-9_z�&��6�՟OjZZn�2�*ͦ�1%���F�p���^G���Z]�\E�1H}ϫ�ciLm��'|�^}��8�꽗�4�?ACZ7c�/������0��onҘ��eLe�1)���]I�6�v~��jc*b-�=��8���-�ɽy=�|���-��Q�C7%4�t�ѢwP;��\pA\��&�.��>LNt�	���l�jKW��]\����V1�iLQ��a9]�f�+��Ho=�ٰ�y�^�j�����}�9�
M�i��Ө�,��a������1�1��f7�u$���!E�l�O��o�Ne��p�o'�l�}r[瞝�s���U��ތQ�*�Ӕ�%�u2�3�(\\�p�B����HD�0�m%�m��b���&3�;�OL*�Sd������h�1>�})����0|�&;c;���!lm6������M�śyj,	�u��}��IM�]�FU]6m6��ű}�j�N�d�����ޜ��}N�Z���d��������S�6�vs��b�41i��z���UKU93Y�G9Ǻ��Ni�B���͆��SL[Lw������I�!�vl�Lj��F����)_{�rƘ�6���0�UU�]2\ՙR�mB�'���6�q���	8��[���A��oS�f����1�F�혯����0��b���ϲ{�w˧��m�q�<�m3%�'�B��뷩$���6���l�ɧ]ߔF>IC[5������K���ILo�b'���1�I,���.4�Adv��޾��r��}z8��Ɏӷ|�4ű��S�ݻ�.I��f��i��%���$�}��=��%�����g1�L_�{��#iN�i#�ޛ�1�q�Νs6K2����S=�.ҮuW�7b9ɂ�����%�1I�}�Ii�QK���c�ێG�ǥ+�9��X>b��󲤣��<^Z�ǧ<�N���ܙ��[��i��v�H,�~�>�nL�$��Bfd�	�E��1�S���A�K�ٯT�֛_m����"�bO���b�~&�C�"q���߱�gl���'��}��;�}�
b�u�8��ݡ(���tƘ��O}����M�9|9��&%�{3��j����z���f�6���0��f�0bR٦3�qH}p��i#�m���1�4�lo��ClK9=��|�}�R:X�hXf�k�#���������kv�Ť�ش�s���L��Z�5)�5��N��Zs=����[wٳ���r�u
����!�"O�$h 1;�����Ӷ7�;�״�TիW���É�%��g���XbY��[���;�צ%1�;�b��͔�쑉�s�&�s����y+�IIN2�����r��;$I��O=?g{a�-4��1v�Y�l[F�{��-"�N��A�1�-��|�F�cHX��:
E/0�j4fLF��ڀ���X����j�����{u��m��!b3z�L|jX�*a���t��`�g�96&�^�l�����$�pq������'�b�Q���c��j��2r���ړ�k��f>��1i1��	lĈ�C�dN�5wH]�J�K|�1�+�D�	}|�M��clEv��U,�v*V�E�afФ�M�����ҝ���e�ݾB�{�,�Lb�����{�������6��s�d�}}~Q����h�B�b[X�S���z���v��G��>�����;��}$��ۭ-��i�o�ZP����Rm�by���;�ILm#�E�~ٯ�,�����8����se鍰k�ce�}uweM3SysWW�����Ոi�\�}&�ga30q�����q�cZ���͘�"w!l}����nI���D��1I����U�18UVXmci~��f���L��l��s�=��52%:J�4X��J�o�p���4�!��~�J�Rܷܶ6��lLA�=���.bD�v��ƒ>v����zr ���N}���imm'���y�uڽ6K�[1�;���AI����_b!l�Y�&�j����\��%5��C�1��gGLb%��9�M�m-��Lgd�>�~��N� ����sf���.���m���du�!�vF
��舡��u"�k�~�߬wW�cu�Lդ]��=}��{?v��+v!�n^{j���mP�)k�͂�K1`6�+3�YX�b6���/A����D�C�`����d2X����2��M���N�v7FR�9�c0e��Y�7�Ÿ٧^�����g�K�o'c\��;�G�dUnF#7�Ym�d�Y�=:��7��l�ڐ=:e6�(�D8U�}[ʌ�B��\fao�������Ct�!(�p"+#��;KM����}��^1�j�'���t�������ֺ�cT�8;>�fw���[��/BM�ٕ����T��${��l��7=�{Ӽ��%�����!�7��zu��-��9�Y�Hw�����/)-��m�-18��W3��M�U�N�*���ަnc�]��zl�z3?Y� S��n>��.��>�fDN��N�1;��pq��q<w=��s�~���n����9��Z���we��v�m-�+���H���̱������i8��I�g�Ұc��u��̝&��m�f\�q�q�*�r�.���5�knB���ZO���!�#�e�^JŤ}���>�clG����F�KIj��WnFn٫���r8�bӿz�;Jco��0[ˍ����^n5�ƚ.f�{6`�`��fIo��8��B�sl�������b�|�i�ue�Al�3��xw3�lݷD����EZ��|�v����Y]0�{�&?'���7t$ZNHcO9��%����6v�����x셤�,u3ڬH�}Se����K6%��U�Y�
C�LbJV{�q����J�e-��S�$��ﱱY���+�dWfTl�~�*��r>9=��
�#�DW��UsS�<�g�=�ٕ�W�?%'V�k>�j'^��dE"��IH��Q��2ۍd��j	T��Ԙ�ZE�`���3�҇��H������m�	t틢O���Jt�IC�k������N1,N���i�6�T�&����̎$o���w:�0��i�m�ݭ!���l�y�N�G�����ת"�13��Xq6��T-������Mu���r1Lm�f�e �,k�r��Hm#�m�1L�H��{_6�&�a��.��$}��q�3>b��>n
m"�u3uhq�Lr�"o�M�tƘ�r�=��:ڼc}�7�m�[�;�onB�hZO;�6�[�Lm�#����ڷ�ݲ왥����1Z�v�]k��L�ֆ��T���{�q��8���(�U$��K��n�4�1�>��dm�nK`�g[4���bӜ��Lj�5Z֢ݦ�%�3��6Ƙ�O���-�Kef���	0[����A��ѻ�bnGs����5�M!�ؔ��[}vŰl�涝�<�i�3�dՙ���S���j���f�ݱ��М�>��RIcے��g]���by���{�^���͋q�9F��2z(�Y���+��"�P�ٶ�0���?��R���w��t�R�ۂ.�{S�9�4��l���]���Mq��̀\\��{�strݲ/):k6w�e�3;�qY�Ňb_Y#���C";�"��.2��?w*��Gk��Ӑ����^��nWg��ّ|���	:ּ�q ���i�R������<ߙ���uG�9P�H%����1�Xv Ә�+��DX��Vq�Т�Z�/S�R��r���z�����k<]!ּ�����¥N���a{]7y+s>v��:�^���`׶�:x��z�����ų�C5+r�^�R)���9���u|�¹1�v,w��nu)�yReޑ�5vIR�%.6����m�0��d���K�����^�o(����Z��ЌX8ąe����]O�^_@��r~�[�N�}�C��1<�e�L�� a�.%*�}��F��t�ht���o�]4�[&-�sf ]@��k��;�V;�@ ��v�� O���+�]w��'͍�R�͠' ����$�kpN�1�ng����]�^%Ȟ��U�ݑֹ���-����![Xs|%Ό|:�U���{;�`=�M�d���^�F���d�Μa�q:죴��ML1p�����̌�͛�u
W�dn���G��I����"�iU�e{��f~Sí��|T9�^� ��s^�dL���jyR�CRI����HW����(�-��(��9��P��n��AU�]z��@ )���������F��V�f�ET�Z�*GE�F�Rv�2��7����LAD24�B-܈)>O��%]�t)[Dk˶>԰�D>ݍ�uB�%i�OC��SRV�
 p9�d��ꋣ��P�[3gN��76)FB7r>I�z���|D�e�[�x��W��,a]�eFxb7#�[Y{�qAz�k����~m��PL;�p|�l'�h�E6T�W�꒥�q���dU�Vx�7;1�x�m�|(0���Vv�jMgE�z�ʬXM�g&U�\���z�ըP��Sk涹}�+4�٘ح�jѳ(��<��I��@ve��񻻍܄R���l?� �a��Ve:�V�	�����u��|�CH��t���t蠙���o����tw�V�p�+6�v�]��|�7��'f�M�6`��hea�7N���[��p:�ɻ�U�]0#*`�-̘��
���E�ȍ(�(�Bdo ��&^�6d1���Ȕ����3�k>���d����r�:IVJCռ+>1�d/��o&S*�O�&<=�}�ug>�**AhJ)�5���6�m)w�ӑ�N����;3U^%K����E��~���;�^6q��Z��.6�"w%��w&�!S0i.�a�'�j]I,k�#����}�7 �[P�-T�m�B��Z_��\m��o�;$�P��t毎H���b����i�6�2��4Ű����d�fw�&�fZ�d��i��g�12�\���թ j&]gy�s��t��K��̬��K�#�h}�ɸ�Mjbҷ��3rRRm	�}�q�u6�y�4󚨭��{{/I���lvϲ(��uwU$�U��M�ls�e����>}�M���JR,k\��LS�IS��;<H�[��}W��;��:�F�"�C���k	�2�RAn[j#�a���eY�4Ť�[)�we����[���M��n��~��4�N�6�&%s��8����H�?gi����&ʹ��l����[�(w3�Ɲ�;���w&�!L��.���U�JCi�}��n��v���\��[~#ʺY��ç��$xBb�)p�%�df��η���}���������W��� bF�J�y��cP[0m6��˥�*DJRE��6�<�%~�`���*������1L̆nE	@SlA��cLF��͘�0eȦ��ɓ���Զ�WFG6�!��vp3Ę��h���~'Q���Z���d�6��������-=�p��c�,A.I��M�Œ��D[�
w;\�8�[;�9���%F�Ml��A�J���z2�guci77u8D����k��M�H��VF��LE�o�l�4:�s�;ɤX���׵��m"�lR[+�����A���#D�Ɉ���AϴZa1),B��v�m-�]�l�)s&�����Ci;�3E2�3Hٟ�*��]�j�̫6�$S��WH�䶓﻽�i)r��񝞺�K�li�w�U���SLm$`y���&��6�ۜ�Dϋe���.�ˎ$c�r=�-���&%kz���4�:~�{�ܔ���Д3�eY���#z���׉Ѵ�sZ��i#IL|W~�ʹ�nY�nt�fVDRm6�����;&X�M��j8*vy���ċM�>l۴%6���~��G�"(D1�_^nWq�*�
�����C8��5��O����Ih��Yg�6* �{s�1����ڠ�T�����=݇�ܞ�g:��4l �l4!� �R��gX���p��\&�.t��{	��̶W`{�.�<5żc��;^��q�����ι�
i֙mϱ��q�=��R��*����{78:�횂��S�m��������^��������x�q�n��;��zu��]�M,2��v88�[��R̶.Fړ[�+͟�'?�"A�`/�J�
bMHbb�IƝ1�H��ߑ���4��u�/%M����0�Д�ǩ��	�U�����Y� 6��0��3���v9�Ύ�6ju��v�X=���'{�zmu��sn˛�=X��`/�eY�^�Ĥ1>׻7`۴���k��4��.2&Bn@���c��\����S�߄~�ŶWR��Ξ�is1����m�u�� ��lo/�f�-�1lq��Q�iLm"��Ӧ'7��"'JN��W�e=�@ˆ��{6"���;������=ܸ�m���GR}��LJ��1����KO}�6i�L!�-į��ij�]U734dJN5'��Z9uU�jeHS�9�$�����4�$��g�����R����h��~��p�M1Iç�RV|[SU9S�a�ͱ�f#���4�-"��d���n�[�
cϼ�rwDm)W�Y����M%'g�B�Ӷ}�Y):�߯�'��i}������m��=q��k��	ݝ�&8��3o<���iQ�\�{'��qJ��}��F�il}�wS�K���{~��z�{�{�PRؤ�{-��!l�{��e�Uv�U�V�q#i����E�o��N#���0N;�J�^J,�Ri�J��e(��Ĝ�*�5��yݻ<��W'i��7���+�<�Wx���Jz�h,F�u����䏘3&-�mĊ���Iq��_HK:2�ˬc�v��pE_�T�Ic������t���Zd�'[b�1n�H,c}���O���%�_���[f1Z$�K�ޫ��\�4L����.1'���jN�ݵ53:��n�lZ[߳�tnq��#�]��L[:>��fjc=���Jc��.���RZS��~��Z���]W�S��wF��WܵbeQ�Ji3߽����}�b
i&�����:�������Kv���9$��@�I��� �"4D�c��/�x��I�Ej2��Jƒ���M�.����;�Iv�IC��7B�)4|�{?s�gY�I��3�����Y�j70]��g�Nll��7��l�z�{n�O+l���W8�>��N7��6�LS�ϳ�JO��%��l��Lo{���0�Lm��ߛ��,B؞c�=Se�]d�eY�B�1�ϵ!���Z�G9$*�4���o��}��[�!�km���Kc�k���z�aٛCI,Ra�{D����ʹ�&�A�n1��Z��O��ˏ����w����yܘ���S�}~��Ԫ���[�h(ur�2��� ������{kr�~�\^ަ�����������N���!Z�8n�����+��Jy��>,�'�I���D�
ӓW ���`�99��S�o�&�oIa�N�M@�ĥ0W���rI`����F�lS����ϙ��ĩM��M��Ǭ����[ێ�6���s��"^&ض'����n)����>`u��Ӧ5YDbVp��ZM\U�Z/*ێ$s��^�e}c����/T�Ĵ?��"�BW������5/�����-����3�[D�ڎd�n�Df� K�
����.��ҕ BmR���j�/��R�L{kG^�3'I��$���1Q�g�;̶�-�m;!�U����>�U����P>���ע��ߟ>J�>�:�`��זS>�# �>]u���H��i�T�����*��ʗ^�]��͓�	V�Ƕ�V�UY1BT��J�H�

C32<�݁��Y7�0�_��VK���*�ul\�"���WhA5��<��$�γ$���_fDc�����r���=��D�ѳ�0�,U��9����$�p�'�>a�"I#�X6�x���fi�RD���gI�9��ɫ)<sӧӞ�[�`�`jh�HsRj�Wo&8�ɼ���
EL��	� C���>�%�'Q��IB@E�������J������ |�j���Q˟�ࣸk����3PC�,�<�p<,�!bMQ.՘!�X۞��c�VkN��条(nϣ0���F�i�)��g~~Unݹ�7t-ۧ�ȟ����7�!�-��]�.��Nne�]#2�ī�W��VH�̜�S���Q�k��Qf�ܦ�q�G�]��N�Ԁ�v��S" -���<�\\9�o����&�6��܄ }J�&�;��wW�&=<!/@d��/��8!bb 	�]Ɨw��~�_���DX��ʺ{>���/-��H�87��m@~�ڭ�7���<���L�3L��+L�33F�q!��Lc�𙥟-�u��f0eWz��[_��	S�J�S\뵟7��s���yh���kV@���3���)�D�I��QbtD�Hk��HHd2R�p�< ��{���t�u����8�t�vk��l�g���<�j��y�G#��n��lk��'UX
���� I�^��ԧ2�VV+��3�5�t�X��͍/	��2�y71��`�c&�\��n��] %��si��bA����4Ek��j�o7�]q[����J?gA���h�&�Y�~��]S��z�9!�m���L���6\�p�y?(J�=����"p�<�z&￰�`��Y3�Hn�\B���2ٴ�0ݠ.�l�2�`O�u:�-�AFMPR�9������ѭ�����W���˗R{����c��ωy�Nh3�(�P�.!��(�83�W��}��>Qq�O������t���'SH7٪����\N��\J���^i�dSI��x����J���J~���P ����.���ua[�x�؆�Q��X�u����M
to˽n�
�~�)>������L�j�?W's'{�&m�a�w�U_Iʋ��ء{y��~K�ٓP�3���������� ��SX�h��4�Î [͍��j�6C@+v�w��zy�_)�$\	eʭ��Y)�t�綔�i}a��K��x��z��Lx�(*�M���$�": �����neo�W}��
�R�>�)�b$�&̎q��\$z{�013�a���:ӛ��m#���9��Uu1��|��y�3t��<��1L�1[����&j����\�X��\���d�~��#��>ԅ'�<�=0ެ�'JǓ,�'�z�Dzڳ���/���>��l��ª7}�'��W�je�؂�c9��q�t^�_�B������+=v'!b��黋V���3��.-�ua���	BU�������萳��B��K/;�/�P}��>?�^SuA�w�R�m�	��awz�M&nA����uy���Jb�T�(|��T؈�-�h?+� T�J��JV%�L�A�ˡF1���7Lٳ\��C��7�aAQR��%�X�M<����概O�Z1\BO���+�-ڻ6m{�;�2�4YWn֏OO���<=
�b��K�<n�����n�\���b��"N����k���¼�
	P��j�3�\.l9:�ٽ�|v�}�(��~��� �C�M�u{�y??H��[�˗Gm�ާ�`����OI���
=��a�!�*�q%��'h\ɼ���U�Lq%�B�s�&'�ZȨsu�m��<��
�[�wt�6~��	�=iA��h�M�D+0_>SN��=��K�S��)ɹ�����K�8|p�ϊ�Pn�VOu(����M����!F�<&(=/���}vX/I�=AH�	6n�B���w��aDG��^z�Fn�Kvkx?�Os���>s�~�f�
�]��鸲ֳoJn4I�\�����Q���l��Rom{�6����_��x��Y��Ļ�s �ꃣ9�$�J hAMWC�C��~��h�nuPMMM�zU��a��5v������GIYO�YL�Ll��+ϼ��;$�u�1p�(��6�	�S�Ԛ�y]]��9�-�T�!r���LM��7'q���w�خ�i�������m�!]7E�5�B�h���y�����똺xj R�Ѝը��S����8*IO\�ߪ��i��U#�@����m���g��j����̫m���Nl���.g4}T��N��0nf�I���Є�$8�0�Y׺�:�9���ZO�$0u��d�I��L3�$������[	t�����V�8H����ߤ���ԅ�ң�Ə<��0u��Z�4�I0�	0�a;�"MA�	��Ct%ʩb�q볧'k�+�bێ^ꘅ��8��bl�.(0��=�p�,���f}���s��'����r����①up�q�z%��I�5" p� �P��_J�<��1�ͦ�2��Z���z�,�~^�u�Š�@l8L�����;�3ط>�!�^�U4���g$���+WpD8�>���U�v���c�0���.(ҳ����o�4���|=���jv{�1�6��9U�x���bm��M���y&/Ԧo�Q�O+��l�	�wr=z[��stv�����M�,ZNp�����=������E�I�Db�Czb��Ș���z�9����-ת������g����Ͱ(��'l���o+p��.�\��#�.�띫#�zg�P��Z�M���#K���
�(]U�g�8�"��;#-��U�l=���Šu!.E�]ݍ8�Qe^��H\�L�n.{R�'��`�0�wJ��ͥ�'����CCצl�`xRJgҗ��}��R��:ܐ���2��t�V�S�پ�02N�ɝttsq;	�Зom�h�vlU�ײ�Ϳu1�N&âu��R�=Y�r^>=���p^��,�Osv)�r|M�:����un^����(AE"�bwtf�R�%��WKVĥ� �9Bys}�_��eL�M��h�Y�u��NCf�]PD�x���)1R(��8����<[�|%*˼t7
�Ι&�����os��ͱĬA��=Z�h>�ն��M�%�n���������u.n��6���╝jc��5�;���j?�>�|�Y�1�G6���'SB�����٢4҉��aKp��Å�Q�Q�{�1�q�?[ԑ?+��l��r�iIz��ݘ���Ѕ��tEeE0=���n��ݮܥ�>=�����S�+�0c�$�/��/F:]��J�q�t"a�3t������A�7���T�b�����N�8��<r<t���s�vp������B�+�2^��v�t��g��^7<�\8�fz�eh�d�Ӵ���1�%J�:�
��6�ER��A�5f,�4eᢒŰ5������v�F�E�8�A��}�pg�ƴkX��th�
ew�S���]F��0CT�rl޶���ܞ�[0J4�3&�n�ja�$�]�v�	�4���=Wd|��i�ú���L�ٸ�f��u��2m��*����h�zm�QI��l��^5��*�̫ґ]��|�Pu�g����X�E�=Mb�$���[�k�q�3��`ԝ��\g��cQ��6N6{���8�)���jh�d��\\s��]Y׍ʊck��e�#]��j�ӭ�k'n�=st�/S��k�ܛoH���+ƍ5d��5��5��xV0*[�!f���8���1l�G���ΡΧi<���dg�nu�5v(��n%�gJ�+v��3A���/�1��8��^���8�7'Z�3����|ѷ��d�Wb�CN��#,��W-糲�	a(��W3�au��o[N��85��ldax3��^���GC����֐�ΡwA���u��\�U9!x=�+���Hh�rv�6�Pԋ��Q���zXC^5z;mS��Ok�]���Clϩ6�]���Z�am&���>�7Nq%�F��f#[�гU�Е��X������s�y�VNx�Rɦ�v�/7�\�-!2��7�II�^b�&�B��r���	�tB��]���×W��kqr�z�i2�2nj��m�V9^ݴ=��3A������\��8���\�᱓g�'Z�v�X���iW��)��8���`#�Dc3�ȸ���S<�DT��w%�M��KD�(�"�j*wN�;�p�W�~�Jn�L0��<=eN{���z�]�u�ai_��C7Z�s˾z�u1AEaYp
girіW$�1�](w��^�����u��,ZIV��><OR��`a���:�z�F�m18�`�D�&Ks�i�n
�U� K��YI.�{u�63�����P��^��WA�n6F��֛��4)�d,���8�Y�!R�J��i�᯴O��%va��$���Է�zw��9A}�SWQf�U�R	iq������p�Ϩ���v�R!�0���h�����B������:жн��շ�>��n3:Āl�a�ұH�ݝ��v��x\HM��ח���R�|�l�;����hb�oM-յ�
�/�+bk�\�@f��t�O�l':��aN]���4͢��Ԇ�f�)T�GoUm�q�+���Ւ��?Z�(�[��u�xu�}�2��Z�d�L�,W�o"�靗Nk��1n�M�-D5D�Xc��w����p�Xl�JqP�Da��!fٰq�&D��p�9C&;=mM/�p�Cc����)@�y��<Q6w�ZGE�1�wS�M���ۚ�]%.��� MH�x��pGC0�V�ه.Vn[�۹�2�$���֧YNݧ$a���t��.=,ƪ�Gnѻ �*��[bzw	Ɯb��nՠ�,��u,P6.��V}�d�ҝ����%��9w
^��Jx��o���%�ȱ����emN�D���Vz�Y�פs�__}���ϥSu;s@c��#�s^�0�ͺ���(��Y>�r ��4��d���(�E����J����ͯ�T�p�����K=��Ű����E t�i��y>�Wq=����$�SsD�����k�s���&�8�;@��x�nlB�R�'���0�fr�؈�zg�R}�9Vg��Uq�q�>��dBN�4[�w5�Q#�`y����������Y�z}�w6��� �(Y��B9�fB�����0�b$��f,>�E8�^'�B������b�;��&�'��EYt���6'���V�Xi��ʲ�-M�i�m#�2��㲝N�6�[���|^��8Ͱ�m۾���v��30/4Ӛ`�o)�c��6���S��F��`lr2�$5(9�Y�tĞ��+�n`v�����!#�L8dG���S��ۄ#�$U�OMZ
\PtcѮb��˥ȠHq�֌u84*��eR:��$������rW$�Z $����;	��4p�&&`��٧c��DNd�!(KELu��>���>�ػj2}Ԧ�cs�>���O�،ρ,luBI�2�	ua����sp���j��Lъ��Ѷ;�Ʀnh7�ةE@��@���MB���̭�fE���[�Kz��h��Nj�uD���r�=#�l@h2h�������ّbK�+�=� ���C}���/.���^����i����H�IAPm�NsT��&��5<�{LRN0�4�����V^,e8P�$1p�Bl��R�3*s�d�h�x>�@�*�ľJKf�󈰨l4<�0 [)EG+g��/2+�oѶ_�:����ؼ0�,`V��3� <���x���$���n�0��	�4�v�t�b��Ҧ��&�ߤfR�Kv��#�/��^=3i�B���PwI�v��6ּ�B;+��0�lg�-Gr��Ϫ�*����d�w$Q�;TS&��f݌i68�D��������R��J��M�p�[IN��T
� G" @"	7��7٪�E+hi��JB *m���뛁,߫�����J��y�N�@�"K���iôw�ن�&�&�e%���$*��p6���;�9�z}Ԭձ�u���J><������)�~�P��[���Ք��8�k���NH��m��mgϒ�by�ǁltʓS!Y{�W���|��ǽ����"�܄$;�&�T�3��!�	"��ٺ��J���j"��f���@(�g���0���i��s
�u�F&�B-�p�S���Ւ�w �#�}Q,Z�;y��x��{�a�v����닻B7�1�CA�!��w��\B�5Uv�Eu�s��Mw�s�y|=�Q��,#�2�iAAc�1�\�`����h��j�2[�ꋪ4Q���}Q���3�7��e����m������=��#��"?|Q����z��p"�� B�*�E���x ��'�̟Re���秓z�Q�� ���"�ބ؄S��\&��G?x���ǳz�`��s�C���A��z�W3�Ǉ��G�D�/a]��]���!�nA�lLl�%�������z��m	6!je8������R1��Q$A�����+�[��P�ئ�����- Q ������{�������"tF��&*�����>���$GQ����u�l��-K5�0/>��Q���Vϳ�ZLa�꨿��}ު�&��}�L4��e�1hxvpI��v���U�ѯ=�Tj9t�p%�Tpň��r�ž�(&��h��%w0=���6��&/���Q�/i�8qTWGӊ��兆����*@��>��E;G�yu�[�Wț�z��i����n�z�˕y��� �lt8oc��&��`����d�M&�l�Bl�ذ.��d�r�ٮݎ��x�m3��`�J-�%��r����#u�(|���,�lQZzk�ѓ���,�]��m�;��nv`p`靪��E��ie�clp�b�]-�Y�-��ڻvL�8�x^x::WL���O/[�>��\p-��ʂK.ᒖ4��S��m��Y⧁�ό���x��G�{t'ä	b�mVN�T�O*cl�˼�\kYAO�4�ً�O<���s�����Cur5��'���k��{]�)il4<�s�=�y�v��&[.�r�i����0"��&.���~��qqV������`A ���K{�?_��1V����׵�(�j���щ#|�.�&�󃈜B �i�wf0��SQ���_��)�Gk��ʏeS����%AJQUV"�y?^g�DA��t�,�F�oS��#�tTM�o�Jn, ׀� G�}�T�˽��E��I/���@��S�a��7ӡ�&��`�+�JH��& ,6��+j�f�����h��*<n��68Z�'�a�{�yf�@���E´=�_TB��*j>�늋a�J @5-m��M$3�иD&�BE�Vl�{ʍE� T>�RZ<�srg���v�SջxU�{�9	�H^ڍ�]s���F�Yb�ٚ&9W������2BI�e��m�z�4ƙJ0�ZS"|�N�2Ӫ��%1�}4K&�&m��*j�fM�#�1�O����D�����5K}�1DX�=�f�YP
ɐ���|�m�Z��L���{޸�X��7Ubm�.@k�U�{�Q3D���HEpf����Uq�u� �o��b�"b���fb�g�]ѝ?4lD��nO
����䁀� �i]	����f�'�m�[�3��^>�}E{��TG\z:8�f�̚A:y�I�q�vu#u�k,ۮ#,ˁcn��j�&�j����R S%&	h���U&�v�p������#�^N*��O�7��V��z � M�~B918h	�5�US7��B�6��y�U$v��ߏS�77�v#�vK��&�f���4Q�K�+u�ȿ|p���0tX��<�᱕~q�G)�������1�@�P���4�����k|�ԯ�d�]��}7��t�,V�'&�P�1hW2��ٕ?ab�ܺ�LE:۬.6�&?2�����*�F���$m�T�@Ԧg��z�ŏ<k�E
d8ݏ��l�%$�b����,�LR�� �限}�I���q]y1B9O���.M���Ey��+w���ϗ��U�u=�o��D��
`��rO��<&J>�G�Z���;O��2byP�2s6\�]i���n9v��|;��U�I��r��h[�
�g��}jνqi�I���g�o�nޏ�}id�UH(ѥ��P=�{�W�Zk���4�[�)�����>����3o���B�`���dv�������!0�F��UyO��A^��i��dh��L�
Iڶ��1��FY��֪�/{�ᙘǽ�%S��L=5��2	ت��A
t��x!�&H��I �v�}�ݕ�;�/���%K��Z�j��i���Q�$F��U%L��ZiƳ(�X���_nC`]�`!��0�ja|��vR��2޴�R=�ADT�3�{7���ޙ�=XN
\��������Jk�Fem��@��Z��Z�5A�j�����zTO�*�	�ȫl9�k��ya�mV��wV�"�=?д��(�!�lU���T�DR{�Rb��Q1D�B!�}�EP�^��L0�0�$�b�y�� p�q��S�2E�;�*(Y+��LW��)Y ����0K,�ALۛ��TUD���/*;��qX�7�0z�=�Ճ�b=#�זZ�*�٩޶%�N��ob�����]�-{��A4�wL�O��N�;����Br������P�R!�BFr-{�� I��ٙD��K�^��D��w\:��:��P�bf��v;��B2�l2Ƃ���V�ʃU�ߍ���` {MW�+t�ټ��WE���q"UF�S]c��Zl��#tE�#	��a�ɊKF��s�۪�;���\��y��2�j9�yij��Qi���`��RI�5`�q+�#Q�M-ا�a����÷GY7�Q��{>Gَ�\���<k�4����F�V�q�V����j�!�I�k��S����-����v�y����%�Ho*�`˒�ɠ�p$">6b���Rl!�$�aa�1%�Dƾ�,��.��T�i�9ͯŗ�a���=b̗���3�N��.Uq�]F\�nA�w���]�V�H7�%����P3ޗ&���>[��p�7���4��j(� ��H�L�m)������>��$��B���޺��6s}S"��>�������O׹YpE"�@��lUZ�Ox�\%��G�p�G"���l�3��J��q��i�n.�C8��bEE�0��C���4{�N�zbj��e|��Tfz�	�yЩ�Ls�:	v? ��.�r�U=���q��rb���hr��k(~�7�0��-��,��Pn�8�$�Jn[��7�q���2�]_dn��f��:�o�v���ET[�jB���!W�ݤ�i{��Gw��%��aiN\BQ��x[ɹ>"�=�!���w�#+k�fEՊ��MR�e�8>�Ԭ�������J'��ڻ ��T����FT���f/����m�,��2O�o꾸�J~�)���T`c�fv����%
���(KSr�3_P�`Ѧ�*d�Q�0",A�%]�1P��LS?1���p<�S`�~�c�6pa�Fq����:���ٟG����p>��}e��O{�²�#��<�4�$��Y@�?�����'ꚑޟ
�_s�54.0���_;H.߹�^p�AE7W*�N���C�x��5S��&����RPE���?������8�Fd�0~@(��6��#Ovf�c��]�V�H��L}����c_9L��\|�x�}��sK�ΠU+�/)��0�aLV �W)�plqF���lU��~�	K���w!�>ʧ=a�>[�}>�f<Eb����)Á���,K����S#�DG%�A������9y�Q�r$\\si���L�E1���>�)1w�aET��u��?Mfs�-u-JӃW���%��5R��`E�J�@6�{v��	R����{~G}�*8������R(]��}�}���_�OLꍮn� Ԗ�n����ol^�����_]q���|��cQ����8ɿd��-�:��i�)̛gM�o��-��ܰs��.X@����p]��4n%}�U�/<s�&���N8·���q�kyj��g%�����|�E[u���B��$̓�2�8�rޓ�6i��K�e\��:�ň�ɸ�F�%m���9�B�]��)��ȁ���{�٠���뽷{�::m[�by�7��#`�U�*��\���ȡ���E�<Q�x�ri�������{؀�P���3j�]L����z��xQ�3�>49uыw,ۡ1���a{u�j.���;�w�VQ�e�P�9Æm��k4P�Y+^wr����5K���ʻ2�j�}&��lЦ譾�Ckz�Ț[�V���e2C4�e��0�O5@�J�7�����p��!\��A>�,��\v�n����vi�"b$�-������j�+��6t;25�]�sX�\G8�ŵw��n���ֱ�A�zcU������SE��2IkaO*ENW&;����@�j
�[>�����ʬ�%��xy��ٌ����-P���)���]8��Ê-'���32t A���kR��+�.J�O�<�
=Ż�_��l���[sua��/�̘{�L2Ж��K����A].�`i=��	��)��Yv���L�Z�%���:�/�,gd|N^�����
K&�+� c�a�Y1wP�)�+v��ԹʞA5�w�n]��˥�5�n�ŨzT8Lmob�8Wm.�~[��Ĥ'D�m�A��)���z?���H$����5�&pf�/�yc�9ݗ찯¼���Z������|�th�wڊ$ԛ�����}�+��謑.�ApjaM�H�Ӹ0	I��CqV�E�F�<a*]tb����'eh���ؽ7��M��!iLcΉ�U�剣�^�K�-��3��Gk­D�6�oR���?mh���	������3�۽J�[�S+�{:��ĻH���n�q0����^l�D�Sܷ.0�q0-6�{�(A�N�#%�R]Z�u=���hA8	~Om���]�s�Ǘ��%�g�F����WD��2�=}�Z��$�J��u�k�}��*�4Xn�3,R�����8ȧ0��|3�X�%r��B����"ll����V�&b��I�O�������RM�Q3"Z
JKwS�ɍ�U'�W�]?2���K��HUu$!��w���7s��.`0�5o�Y@�$�V��6yP�{�QTqw����1ƌDͨ��> Y~��k}��\ �N8`���ޯ�G�>�����UZ�N,�Z���_���X��_�ϵ���Q����{l��v���jjk��wi�ff�'������[R��#UpV{�14�C�f����S��gՑ(�`��w}\*.��;�9@�%���ʅm�W_��/{��(@F�T��it*�oM��U��xo6x82�F��w��]V]��bɅ�NO��qmy���9�5Tno[P	�	��l�X�|>=1@�]Q��g�f�J(s�H�k���oo�d*��^bi�� ���Q_-Ɣ���X�R�eV�:�B[W�;��ˏN�
��h��/���1潲�q�YϨuu�˃�&��W�/�*3C>��LC��Uq�EV��[�M;c2{�S�
b�T����m �`��U�=�k|zo��C>ͅ3�]���q���K��~�}�+�*&JKJˡI��-є8n��nJ�m�/0��|�n�'.�Rz�|��bTZ
��-��^[&}�S�Y��}��#@l*�uF�7Ǡ�l�Y��	]+;��S��vOEj>�LҘϩn��d��ը���>͜��2c4&!&a��i]_���&�&Ͻ�`T <v�6�C7O�f2�y����qi��	8e��f=�/8F�%�����K��bi����E*.��ި�������*l"��!6J����^�7�F�^�������#T1~�8��F�We2:R>��i��J�1*|#1�<qh���d��THޥ
R�ڍP���B\�?<�+6���:y6c�d�n�8?3�F m�j&�mÎ��j�kqn��n����	f����V�љd�l�qc@cg��l]	uw&���m��y�,QH��t>��]���B��2�eΏ�8'jI����:��ݝ����q]]�C� �3�:	.�jه]\�i��*�N�St�k��Y5�-�,m.3�=~��'��/�4Ƈ�i1
}������ӕ9�ӽ�ϮL�2�c�ڦ�1N�%�����|���N��zpB��b��'��w�\=�NP�����h1�.�t0�y|���춚" ��!^z��h���2�/o���K�lo�6*����<�
|��Cb��O�i��X�8f:jj�=t���P�Q�U{p`�V���$Z`��6�L��>�E��Q(���?z���VEK�J����O(p�A� ܲ�5|�@"��=f��}�hR;��3W7c/;@�y��Eb#�r �D�wl^��*h �\�da��Ď�sftʥ�[4��o��9����~{��hjV�p�ぷ&�W9���WhZ*�F�����"���SE$l4�g��IUb�O�n��{�Bh o;_*��R�bЫƪ�%�a:�p
���:"��M���m�nLoZ�j��4���#!�/G@�t����U��1��{'l/(�ngm.t闛�K6��"i/��T�*��);S.ߒR��
`�=e(Zw��q�Zi	�s*�wRN�0���DQ(U��p ��%�U1J���w~�>�������O\r@%�J6J.���s�1�W/�µ�3��u����A�Q���� &Z��g=��uq����j�Ӿ7f�ޚ;~�P�dHʹ���ø Ai��PqTA�y>�hG�[7+o �^8�w-�F����j�$tϬ�֜B
��)�C��'�بa�IM�m-!\��WR:z��cЧ�/�L��`���;�}R�Z�UW���}� Ǆd�~S4�w��I-"�H����k��=�<>1�z���@W�"��!�����骇:�P��9#�y��6
J�\.�QTM�-�0�e�"�L�ʮ�Ү��JL��+%��Jw�;pǷ<��	�����ݻ�+\��s�pD�f��|�z:������8�q�L�c5Mc䵩�%�Tѻ���IT>c�܆��u��)�־��:�?]�gʕ湣Fvt��C,?�D��f��>B6�j.��oW���Ǧ��Qk���\P�
�]��ޘrv5��$�%�B!��ص�/ƕ%	У��ɯv�N��g|j��< �Ǵ�@�� (��ÐNz�ӭ�Q��U���k@��vl��M�'��=w���G�
��*En�\���ήT���Hoʠ�W�.�*K#D���"QwH\����?w�8�$iQT���\`�����)FڏnA
�\f�R9�a@I�U�o�U}J�k�����u��@�{Fv�u��Y���7'	��݀"DǏ����I��!����j�j�k��3o�h;��v$�b>J;t��vj''=u킫��fy��A�e�dǑ,��y�_EͥBm�X���aެ�m��!��X��k��SV���m�[N�c���Ǥ���xc����0�Ɔ)�"T�ܙ;�����]	Lm	W��e�U#�iP-��-1'���sFx��o�a1�b;�q3k=>�Qpm��Vզ>��Qڝ#���a0"Z(��%;o7Z566�'z�G+v�7�C�n��-����¨��T:�%�'n*���@�?$g�Ӫ���2�'�QEEU+�x��D�P<mʓG7]I�~�1[ P�V>��*(!(��RY��3 ��3v�}��;��ެ��;�t����\j�D2����1��q���}{��K^�oܪ+�C&(7�&8��ze�5I�ϡA���&�,������/��/dW^zMP8{ީ��gL�	�"��Q���G�Lzz��C���}3��L1�:�]k�:K��X;c����[8w�R��p{ϺyS�X��5a����`����A&�/M���Ce�`�y�K��2�bK,՛Yu]���AN��A��5�;��[HY���S���dI��V\�4��Pۂ+�Kuܺ(]�K�\R1��狈ݕ�Y��&�<��ek
�r'4R��x:��9�;�v��r.nnx�L7Y�1�&h���<���i�?{d���ƀ����x�'S���iM�,*�lbj�Yu<$;L�	1�.�[%% ˖�dG}���]�8@�9��g��`��9y-��>����,"� �LW�n�D�R�S��!���,KB�O�P⪚��7�2X)4�L�Z�S�����"I�]&��������\N���M�RI@2	l�l��^��T!]�QS���8����.��z���Q���Z�ZEn��	0����OgLURĽ��uT����D��f�k��n(0�iDڸoz��ujc호��֑]���GTL
4�x?w��h�~����������םײ���U��a�砜�;�e�;0��kM�|��G�w�j)g.�T��j=^�Mƕs�=f��G���XPӄT1�uhﺀ��.���\�|� �K�_K�Wt/h�.Ki]7��-��o�ÇEצHcoʻ�P6�c��y��4��ڳ}W�ns�P'��K~��(  ��?��􏤤&{yG>uQY'�K,i
t���
O��$wy��"��HS���F3�ҩ�������5b���d�G .�|��ZIa���oTUR�3����m�;���x��˵ੂw4���yW��&��خ����Q�4j-�Ɋ�]��4�����'�:��qyH���ɲ�5-$�q��~��^
ҡB1l�Us�.��y�*��������Ϯ��쳑��ψ�K۵��s]��Z��ŶU���/���jń� �-�X������ԷܸW����r�v_��kN��C�YH�n����o��@t@���&l"��.&i�jY]�8t�� |Qb
h�ߗңzk�}�wޛ
nc�B�󬰳MjL7�tP�Teэ�v� ��SF�$�b[�oF����tf��Uyӳ�5��+��+�)NgQ�M0�I6t�������pVc���~z��[8���M'Ë���}9��P�����"U��s�V�:���Nyo��T�<�N��	��6���7.,sW�ȥ�i�+�*������c*+�6=��������na�iZ�@��4��h����N�h��߿:m����|m���Ow�~���,��p�q�k0�N��������uyf�4���~G�7cj[�#,�s�Yú�/k[>�Z���>��yF��94c��pɀ��
�S1wAg�QU«�VD�+�7` ������F��%*�q���
�U�`�	$����ަ�e����|5v���s���*a����L���&Y�3�}�����U�C��4���w��i�[��6�r��&=w��VGF(��/���E��x�
�c������@K���U���b�D��z�<NY�2�CF=�[KH��I��c��bcJ��K�!Y����E	Ł�5&�m���c��JH&B)f}6{g¶����>�g�9�g:}DU-Y�[t@Q9��Df������[�r^QM��JM(�!5�͑���6�8Z�dna�ˢM���j2������Z�T��� ǆ��o	'!���~v;o��:(�����Q���N{ڡ0G�>�ulЊ	"���ꊑD-�ꕔ~���g{�Id�N�{��y{���}������LP ��]Q�C}�CԬ��:�n�TMU��Q�c�Eϻ�&h!���vl�z�E\y{�|�,ױI�t�	��k��l�MR���w�
�}�6-���wJ�}Q5T��E����Ǳ��~�;&&��F&tmA[�Ů�1:s]['`���]�sa�/`��5�-P�O%p�\��%�!VL�\ND��H�2q��N�I�X.����Lb�whG].U�[ΐr�ɝ��r��� �T���mph��}�uupS���3l�yU��|�bV��Q�7|.u��O�U��nphMz�z��7.w+;%��g���e'������m�����F���5�޻�2����^�-��9m7K���p��N�)ZWf�v���/�U�QY,PcB�w����_q2r�34�M���Z��W����u=p&o-�u���������;�J�&�/B]F�8����Q؜�[7:���Г��6n���Q*6����ք� ���3��01��ǰ��n�H�9�rc'�\��,�&��y�hbU�/�2z��񮐙S����\��z+}��^�N���͡�U���X�:y[�>��d�,��Quu$�
�;��EmAt�ңWg,���oK6F���2!�q<3KږM�AT-�#~�$�fiD��45��*��Zb�R�j-j�d��sEL�4�z�F�fSZ0L�m�ncr�[�&�mi��ye�pQ)lY����H�{x�?J���>�D��r�u�xY7����Y�^0,����O2`Ij�xf�6�?u�^.�l����ݴA�n��~.R`��n�}��6�ǥ��fЋ��wK�t�rz���[���c�ۭ�ݲ�]�-e�����Ƶ�&1&��Ӯĳ�1�Y[���G��.��F&���T���ⷵܣ�s!��S����v0���q��ɇǆ�d�$ueSX��ZD,,�`bڣ�Fӧ�Z��8�3ۖ�K�q]���l���`z��bQ�x뮫�AƼ����닓ns�^����K��K� ��Te���cr��u�ֺ;J��ܮxMV�T�g��R�	�97m�Ms��ٶ��nM]\��(���.�V�p�◧U�I����役67i�m����S�4��E92��p�-��NټwGZ��X)Z���8��5��S�#y���r>Cf���^gɪ���q�s�xH5�tEfĶ�:�`�\����Z�Sn�ZW�����/+,�:�p爎%��s,n������:���i���/jZ�;u�=�^�v��ٌ9v�bK+iD%�l)S/<C�8�\۶���v-2�,Z����F6�J0�b�f+��i����i�kse��ҲT&F��pKk0�6g.����i���h�0�7���Q@9UMۇODW���m���烛l�rխ�緛s����b�T��N{y�Ǳ��@-ڄ�G��e厍�PB�lҷ�pܹ�h�6ј;Z�q'�Y�.�=sc<k>��X�d�ڧ��źx�w	ZGz���Okk���\���{m�Q��G��GEƤ�A�e��zc�W��\��ė;�C�`s�Ox�7g�jv�ɣ�5���[�β�K3L3]`Ig�Qmy��I������m���g��e������k�۰�p弮gR��0����=/eł'S�R� A0	@���F��(�kˊ��B�K�b�
��r�e`�g7�����o;Y=��U�1ƒ����uh����k��rVs�]v�w���������'~�|����xp�34]%Z@�sw��`��դ��0����R�5Ψ2q�62��*����+5t!����^��v�eY�O�ǽ�v
�F{]4�O�1|�;�����&�Ugۓ:�%�9u���ec�<�!�
��G�}�o*|+|�/�9y���mqB����лI�R���H(wÂ&�s�D���ys=����۹�8(+7q.�����g�Y�k|蝸�I	�U:���_e �m��bL�Fw���^Owr�6���M���Y�^�8�t� �~����kV׫�z��u�k��<�cQ�t��mi�T�J^��U0��6����:+��qd�9�#��X��T!l�2`�Z#㼴K�x�LS A��A���={�"�:��Q'��^-���&ee�wp��n�v����x���d�%����3ä(��8$���b�I�$F��*"���*:���VŔ�l6V���O�P]B$���!�+�s��ں�'��T jX��^�0��d������՛p���%
o��n�xZ,<Ҍ� ���3)U�R{��Ď	A2zTÈ/qď��}�1"H�07n�HX`��	�1����(E*�\;�ɨB05[�ro�Ll�4cы�߻��_%���1D��6��-le�Q灺�W<�a�ۙ�勲]��&���t{N�Ⱦ�D{;���cs#W*�+ͼXK�t ���. µ�iyC]a�[q$'�&��,�1&����{.`
ʛ���aݗD���ʂ��2Mf�T�K)5()6i�Vk�5��v�]cF����z���ődJ�xg}%W��\-B��Io�^gN��l�+I�����&9���F��=���2���
=�ۉ�z������e5��$2ݧk�i�l�d�b��[hP�_ َ��.�\Zj��m6j��_����x2M��΂����9$���LE]���2	&�	S��{�~��Sh&�Gzbn����y�!{�Փq�� S*�3�5�,����	;V��q鲂
��a�w��;.d�-9Ɨ��$�nI#�@mC�\]X���
%'�b3���vz�/z��|TrFz|&讎���Z���_�u9"�\��߭�6%&�Sow��\`K������}z>�[��Y�l���"�ժ������FW����0��dK�T8k�Jk���UM�tC}��5�D��wU�E%#��e!���2 �%&��^��)��>(���|��;/wUk�b(/SrNh\R��箳��\yK�f��/!b��vX7���,O�/B=*�_��V��>_�m�q�/ϝ/$�1�I�!��x�=>Ͻ����S<p���g��Dz��漦������:��V}4_ve�� [j�/�z���o�t�.1b#�gE��Q�ޏM+��5T�|d���e��0�n� Y�4\�g��J�YԦ��¦��1�H�{ق&�( O���w���Ve��L���dꩈ�X��>󊓋s�we�}>�T����}�-��0�Gv�%ۛ��q��j�GYB΅�5�p`3�D:��&��p�j���1J�xL���7��@=�ݏX#+n&��W��Ș�@e�\]��O�n�����M1KOw[�s��>� ���"��-ꊁbD4�	�{�T�c�U���ﰖ����Y���Wu���6 H��y
d�[�1�z�qtFt�j��b{U!h��\��Edt��y���H�B5�&+��u�q/�s-I1�?d���1)�L�]�~�L�6��X�#�тR�	hb�Tbw*=TW<�U,.[��8-2�K�N�pX�M���Y��yx7nr�L?�<U� ���$���<�JP�J�&�g�QB��"N�6�UZ�ޚb)ު��םI�O�����:��h��(��+��V��m��5r>޿�x�U80�hɂ��;�4�gd�>�{jqzs5F����~��(� CNi4�Q�ޞ�"Z`��ulԚ�~�G5�N�d�LI3���`	&� �-2,�{��6}�.�1,��*$>�D�J��w�U4�}�WBDa*b��ٳ]�N{�ELRQ�5����G�LxDp��T�d� ���({@M|�\�J5���'�`f����g�=�"+]�F`�'G��Zt���Ԇ$�Ṯ�����{�v�>~M0�����fd�9%\ÀA��! �'��T}ިQ@�	��wϻ���,xznv3�3�׳�"�;�Nb�Ӣ���Ն�J� W���t���5�4�F���í93=;�\�Q��|�� {+e�	2������>�ߜ��d��_vO��C�]]-MU�������H�N��z�$�c�@X���p���5UV?N̪��=Wd�q��l(P�$��ި��E����t}p\`$O�e̋C��Q&�s�$)[�.��C�1����d��*��}$m+9�MӴ~���*�g�=�.�9G�l��-���#����w�LJ���T����0wܪ�nEZ&x��g�^��q'}�z����|��@�K�W?�a��j���"G���.��o��T���>V|�Ԛ��^]k��0�;bJ���Gg����=k�e{��ļ�R�ɸ�;r�v���tr��3� sDk���Ɖ ��m[������3��zmk3O\���6�Hl��`�!ōiK`����^�2�:m3)68�j��L\el�$uF4�"��3YN:��� ��@4�G�"oa�z�Y�3;&��&���QH���@hѵ�F/�<y�"��n����UR96����)�V`a�.;Rgq�u`���:u�@�n�^�KM]��9��&e��]N��O=�^i�wTURy���'|  ��5�搃y�\�e ������ڍX<�MR^׮�o=U�M�l@�u�\M���w,�����ևo��}d�«ϼ^�g�j��/�Cy��R�װ�i���e�����<�=�Gi[Ӣ���Eu(�u���z�V�Z����(���F����$P�7u�63:V�h}�Q3kϧ�B��\J#;��h7�0�Gb<\��Z��9��Y�	N�K�_��G�{{v��O�����̈́<����o������z\�a�/"[�0Bj���q�Jj@�G��ƞ�
̈�۾�7�I.���A8gxa��2yÏ�B��Z[=��(�!A�A��U���r}�S�"��]�s&`�Ƒ�"�'�a�� �bv@�av��:�L��̝\��S�����rh`�<*&� �E���h�ZpXM��ѽ[�]D�B=��ySN�i�qT~C6tT��sPE��qm4jv�%J���t(�Nq����u��B�Pb�}騚J+�ǣ��d$X���=<*b�!��xLvu;�az��7g~��HMy��Uɡ
N���a��$�Q\��Y�׷#�Nŷf�N4�z�wY兙,�����><<!�Im;��>c��s�B�h�4�xf1}\��\7� �FH��%�~{�S���5�%2���w��U%ۼ��F�s3>p^L6 $��hoz\����犭�������E������EG�C�ʠ03��T��m;SMq�B��>>ӎ���uO9'���c�7�\��-�Z��SKZ�O��չX_ф�17yP̃?@)�L��%��bM�1��i�\$�D�u��#�H�q˯�K��uqh�4)
�=��}�'���t�ǡ�i
b���O
�^Q�|(�/31�w�U5>��To����^���	Ed&Ӏ�s�	0ӜY<Lot��5�;P�+/���cT��Q��)��VVo��X���ji�N���©�b�!��)���ɐ<z,K ���&e6w}W�}Ù�˟G���!/gyՂ,��P����ȶ���|�6��`��k��KWi���:���\\Y��Mz;j8�ZKa�uh�y_UR}�X��������Eq���~���|�a0F�j�9�W��� ���v��r���]GWNoq�����7s��*3V-9���7x\�����~ϯ�6Pp����<@��L���u�u�J~w8�x$�R.]N�8@�Z�B&2�k�X��N�E�[ 6��^K�W��¤���A;V.+�������j��:I�}��2�z�1-cL!F�����[u���l/nq*P����q۾a�m���|�[�ޕU�:&�{�
���� z}F�%�w���0XM U�����,@|��\X�`���T(7�[y�ut#"P7�;��
l66�wOޮb)�<���<[�S���rj<���4"��	 Il �I�V,��-�˥
0'wus��׵"io�EUG��p�
�ˣ2j#9��J
i�EKFw��}����Qrm^����4���{��Pe��QU=?.;DG��*��1�����f�!�%)#��B��-g��ّ7��t]�Ǽ�w��E�SL�S46���;Xm��tT���-�&��۠y�*g�rd�j�\��R:1n�a���H�U��Cٷ����r �����#��\�W�������,�w��5ۀ����ea87��@���My����kݬ&����f#�7�����ĝ(��Ivơl�˒m0o�����/Q!�'�31h�B�c��I���D��y���� �ǍQ����[Z������{]��"�UΜ'(k��E;������ѡeD�'�!���)����d��]
F�i�"��j����?U��ďC)|�&i]Z���|6���ǠT�݃�oz��<ͨ�`G�ޙ����p���G�? �&���p��X�D�s>�#����D�Ƈ���B��{�цBp�C%��8| nz�EG�n�׺tL�%�ʪh�y/���e�SMcǒ��R�0YL)K��[�'Q��*a�ܒ�DO{�3F%���!�[����4���8˸���sC��e��ZKV�
�ڂ��^��;|򭦂e�[��7��r��G�m)4�<���۝����T��|y�SH2�(�\X�=��wQ�Pb !\v8�����a
 ��v��(*1""�(K�2�Ҝ���}= ��*�����_��+���D��)*(z������O7d]D�����L��FD,1T�	`���*�� � gS��?q�T߳UV��]+;�t&t�`&HH�32�j�zhTWt蚫Q 8��jώz�ݭ��ѯ�͎*8���W���k�u�S>.�!��СK��!Uj�N)�&�t(�{��A�+�l������'3.m1D]�����⨡^k�� "Rp�,����<��&{>����^'OS��sM5���������~���Z3q`��}FM%��B�<��"�ϴ�U�Qb��c��(-�L��U�}�[��'g#c8�}�%�7��]�sޕP�?H����d/rQ�n*d�u7;=Ʈn�S��H�gz�)1�K�eӺ>��VA�������3�r�Y��ˤ�',��J�a��8^�/�=wzk��:T�ySp�/�U��6�Gg$�tPN������yB��S���{�,���軤ʤa,�2�MZ�\Lu��JCgq�H��깖�t�7;R����/N>Ӵɔi�YW�u	�ME����-�u�B�L,�����;|��˲��2U���ys� �����:V�vw�"��f1�5ʃ&�3kczXp�E�j��_:����6�NA��a�J��_�c�}yެ���\<c8�vK>��%�J�u7Ӡ�׊�x,{��L�R��4vͺ�s�铖�/0b;���G�͇�ҭ�D����D��`�~C�L��ȹqW((��Z��+v/1�k�Vȁ�Q��<���3!:� �VMu|�u*yH���{CR�{f4ze.�u(Y�:G��ĹAcb�	�,h�\V�3��ʹ�u�y%NT嵊�ӹ�Нݛ����iM#u���jI&3��Ո��H�*�hS�u�xV:hv�/�_P�|�!�[���j^,�YHk�,u<?F�e�:��!Z,v�y j��Ț��B']uk���bl�����d�Ҏ��ضUZ����_X�:7���v槔6���eq6�M�#����Q��Z��T�4��
�1��̽#���;5:w0,��x�L
��*�ұ��@V�w2���eNJ��^߄�Ɍ�q|H�K�US���d^6ōM;�=4�h���p�� ��>�j�:=W`��Xp�����C�s�#�� ACf m��;\�Q�OY�|f�v���k�R(FV/�p2���P��&{�owM���N���F���v[��,�9Ԩ�rl��ߓ��p�l� P߱��cD}��>��_�ERmE}V��x�/\�,}�@�X�Od��M���
U�G�"�-�O�i�.� ���ݜ/�z���b�F7���S��Y{=�յ��ٞҀ�����A�r�$F����ɩ�Jr�VR�.�E5�	��G����W�:i�:0Z�t��.�b1�F��ence��M���S�1�>F��H��k�:$��'���i�B��v�@ .U�4��k�VV��9r�����R��di܋�M��1�F�Q1/��`�ҝ�r���Gf�ݟ>�5jܰ�ڧ^wY{��:5kN9�����3��Nח�ٛ"]�\�û�;zV���G�1 �O:���O�\٪�6C�S_���yrK�vگ�˘�,$:��m����V�޶$N��ϯO�5���;�;�CTe'u�Gݰ�>�N&2h�^R��)c�=�-��MZu�r���9�~��r��*ṣ�E�����5o}*�5OP�B��ϲ����ªzW�8����J���=&ӯY�&q�U��`��,u��2c��n[�@��iy�dC������	~`;�m'�E������P4�d_]l�>B&��G@�$d:�A?=T�O��u9����"YM��eI������/"��^�����u9�fnw�u��Fю���s�4n:2xqd�!��M�գ�����Q*fv��Y���>��f5�v�b��1��Ϝb;Uh�Lî�g�5ͤ4�ٺ���K:��|���A��Ҕ/o���yҪ�X���.O1��]b��g�5��9��i2a����z���p_p��h{��+EM�u���+&,oK���������m��n0���!k�yU����"�r�S���2 ���.��G��/p=�$�0_̤n�!���_5PGԏ�ݳ�n=�1�F�y�q���$x���@��B�Y�������Z�{s�ܴϭ7��.檵x�:����O��3����-�<����'��L�P���WG��' Q"����NH2e�Z��!м>ކ�P����7��EX��>���3���Ʀ����I�����2��&��P��Į8��u��];vM̡MSY��e�|훨��F�`�]����QϷ���s���F
5�Nk_��0_̈%�(�vO��k��1G/W�����˅�ޗf��15���]!���8Ĩ��pWȤ�Յ��4��j0���X�������UPB����
�0T�e5j�m^WY����TL�.�U�>C�l�[���Ǩ�� �����EU*���j*q(������״ �-��H���6Ď�67m!D�I�	�����^�	'bj�v�G��U���Fm����v�s�@�읥Phc�T`dO��P���l�n#�]���n��u�k��J��w[�,�&2�h���n,�aU�@e�@��6,kSH�Y��ڞ��'b)�v�$.��֌le�����#�s <��]��<�cUv��s�,��t�5����-�bX���SW1t@�x���$�
1�밲���ſ���|����������B&�K/� *md���7��p���w�v�e�]��CϗמOV���R�Z�m�M����a�A��%V�	�X�ڨ�)�A���a�7W��=>v��w���[DԘ]��R�3&�v��P�`AA���Z��^w��Y��xC�}w.(�w�bf�-���`
�$�:����͸0�h&�!��X����/X�#D����A�ְMU�Oޤ$�}��4n$�MX��<7}n'PN�
�����׽Ψщůӆ27LF�L����wYS��h�Z Ft�T�=�/W���,J�eѯgLL�soO���F�f�,7	�-6;� �Y㛰;����6��߲x��K�6�[����|�I����۲��'G���� n�������$� ��y{}5�*�c��Ҩꐰ��Gb(+3��t��Y�E�"��5F8Юڌ\�3�v�:��q����
���l�q��bE�ӧ��y�vh��/�w�X|Z>��  H����I�(���p�e
&��X>����r����zj�@�d�/L܂	�)�ۻ�+}�UH��U?>1{f���̑��4�=���H	0�]�}z�I2[�򽵞o�����M�~���]r<��I�C�
̕�C=�L�A����H�ޚ~�TUR��ʬ]�(���"lR @>$B�"�j�ci�-..up�]�k�]�1�g2���ye��'������;�3F�q�5�q�����>N��Ԫ#����$�d����QU{��Ǘ3�����]���S}lf��G۹�DA�tn�.���3b.-��qWJ�oUI�=�n�(�K��n��z� ���z]s�}2�埸Ov>X��5�f�x��(��$,n�d�)fn����w����<>&�Q�~"�ǁ�q��jQ2��4�A�i��tK�Ɍ�7t"bo	�72�vJ@� 4ߨ���D�TR�p���Q)C	�n�ｪ%%�2l��3[��5U��&�z2��Ȫ���(�Pa�S[v��{�����4��"�W8���缮�{_��.1�P:=�&Z�B Y�C�p��D�x�qq]�F�]��)j���?_�/��=�^��^
=�:M�f�X�
��Pr
�z��ш��Q�B�����ƽ�̧�+ y�M*H�u;�~f}�G�½�La��#re@-0J���3�T%�n7�]�F<;��̻���bgWz}��ߣ�#̒��Vn.|�eE�����}Ƣ�%^ͨ��W�.p8�k���g���z�P�N�e�b;�K#��g�r!ŀAڨ��r�����wO ��Y\	���3 #��)M����2`�9H}q�l��v��X�1�̐�s.b�T�'��mJ�l!��6� ��J�6c��F�N�x�5��v�Ws��9߳Nk�GS��IݹҢ�f۸b�d��Go7��]�l�������V�_~Ξ��O'��a]�L����bz�d�&�^��A���I�v2�����B.	P�M���<���~ ���>=.����tX�O
�+��1�싻޷hR��A"	kh��]&{'p���$��Q�{:��q�=��ʊ�`!�� )�ջ���q�?�����<Ч�/���F%�qcq3޾tL{}��!3�S��J3g�6*ͤ(_�NEO?M�G��銓C_��o��BB��0d��^C�F'Mc���'t;PoL�ׂ3��&���x$K��cB��)�N����%(�
`:�Z�9�cod�T2���i��p�gtr��ݹ�0(���]I�W����["�9"ŉt{s�q�Yz�J���h��A�5���a��F.�5ґ��MLj�WW����ufy�������Z'��f��g�� �v�shZ��+Xa��l����.��/��U�F��|���� i�Q�Io��u�4�dJ	����>a��`*T�P�z�N�����(�%	���QYη�.���d��f���5������cG{�c7̤'��گV�WM"�۷�e�qS�}�,v4xz�@��bh��ir�z�����d�(6��9	mυQś+�ѻx�v��)\v#�8?20�Wj����Q���򙳳��};�Jyo��Ӟ�߇0�m�@D�s2�k\�9�GJ��GW�)�["}��r���4�쇔Ύi��$����>>��:Ss��}���x[���q>�TNY����&���>c~�����<��z3�姴�Y��y��|�$i�랗��Kw�����B�]�r:�r��)�Ӣ��^ϸ���d��/ҧP��|h��-��+�����ǣ�~�xV�`)o�r�ܟ*��$ǖ�@�wd��y9�_+8ʩ]?�q�p%VS@����8�����~��ѣ"%b��%G�f*��p6�@����p�4����))���
��sH�?m)"�w-�������0p0LN&���~�=�5<���݌����=&��㟴��(��L�n�Əx��ɫߛ�����&k�t?��F��B�&i��U���P-4`�I��Sh{��E�h��}�K��&b�@�oz��G����rhV�i6�3����5�.�rv�I<V�r��G�!_$̅ �\2�	Z��O
4��5�U��O����D<����.}�I� ��	j���
3�l�,�ڪ3���QL�{:�M#���g_�}2�E9�Li��<�@��Mc�q����r1A3�޶��Ho�K�r��t�eh�������e8�/^J�L༊�t��ow�k7�'�~��� @������|L��[�v�i�
64d��1C��`�6�����/d�MQ�"��5�L�[mT8�KO�G����%;Lg���Y��{_�����H^i|��.e�Km"�x�<��uXzb.%y�j�����ϑ��/���*��JD��?�cR�%({Վ�c���4��И��h�R�%l���Om�� +c��d��9]�O{�뱢��3H^l
�:E�n;����_�A�(��a��e�}�W]��ԂM�yЪ͞����Q�Dx�0�S����Aa�f�2���Ts�5N��}�Ȩ�!k�Pi(հ<A)@]�PZN�ق4߈Ʌj�{�Z&���ާ�6-{�澼?d�LO�&rF��-Sa���g�{}>�� �5¦���\���',�C��؋+�a5'f<&a��EXWn��>�/�L!�3�O{�'�LH��,'�2���d��k�\T��MnlI][ ��l�Y�x��I��nRI۾�mf.�~|&No'��7~�<�Xng1�k+bJ9׆��Ѳ)vM�hw^�!���i[g��۳�{�֦��v�y�{zhm!�������`�@����{ƫ�
�(84��z-p%J�7	�Vȋ����>uf������>���A�I$˩�T��m�XEU����ª׷�T!Q����Vt�4m������l(L л�12 }���}�Uv�����s��t���Ț?-��H��i.�-��� ��_�Ӕ�[�*j������3�&	��XB�����<�ɨ��p�9Y5;u%��ἏpJ�z���Pkf��j�j|x�֋�m���5Vqq0Z�PdҊ�ܫ��t,�jg��⛭V�鮳�#Bzo{��T��}O6ߵ�45-����j�²?i׶kg?�G��BE��U�����t{oLQ�kU��Wf���M���JЕH�T�%ɵ��$�����V_ .�]2�ʓ�
z���
��K�y_�L�� �w	���}u�}����Д�J£x�r ���ӻw�؏���j �wT��d�ے�j�K�J��SR�~����PN�2�'�c�v��t��'6��:ץ�2���ˠi��=�[�������,�Ã����h�s�z~�t����P�X{Q�WZ�������=ʗ�TeJW7K���Uj��+L���X��h���P�=6��T�s{dF���"\�ԭpm�`�֞.���]u��x�T�����&�ѥ�ؘܓ��8l*Ó�@́$ꩌ����1Ӊ��3�m<c�����Y�Qc� ����ȭεߛ>��^}����*�5��3mV✴��IѕVRw�fm�k˶	y�-��v���u�}e+N�Żw�ͥ���Ң���=ץ�ux�I�R��K욛����&���w�o�jb;k0���m�2E�������t����O����p��Y�]Ft�ː�u�n/ݵ\킶
|�n�5�[�*�E@�� �ĹtU�	��k��-?�� c�nE.�祺��I'*��V]t±��ܚ��r(���emGizݩ����5<��>yq�̫�����GXȘ㌶c�6Ŭ���C��,;nMuh����'m��ܹ����'s����M�� ��kv;]/a��o�:�dRO'fE�n� �[ciY���tZlq�*�s�
݅�7h��kv*� ��V�[�:���΍)�FՓpV�8�	����f�t�fN�ܝB����k\;4��,e%4mҺ0�ݎ�t�u�$����=��v0�:��B#�m��i�Ogs֥ӻdSc��p�F��-W��F��� �;bN��]G0-��,i{c��zf���9���졮��t�o����`&`�,]lm�6�WK7��ƻ����	�lw< ���k�Xn��#����g��c�n�P���n�]Ev=�qƇD��9thi�kn3r\7j7WS���R:Y�R����SX]!`/���ܛQh獱�Ei" Ѭu�c	Ч[����X<�Ɔ��l�^0�Hy+1�����٫�`�C�؃���Z6u��5s�l6�q�mf��(�<v���3��ḳK�A�5�u�.���_l�6��޸6r��� �<k��[�W7�nu�/ K!˦�V�6fu[0jL)Y���,�w4�,��j��%����Ķi�ce�4��[�ޚT�le�T�(���Ԛ䤣��tK��űBb.��e�^+1u����F�C7e��H&,�-��,��4&�6m�G����k��#s Ѷ�B�.[�u��q�^�j7nܜ�k=m���rM��ҹÛ����TkVT~N	E@�	]��^���(�Nt�]�t��\e���э�%y�r����S%��塒�6�v'"��ʇ��;��R�mۦGf��oq��ཾrܮY���{�6��9����QV�x�=�\˺�]���gu�}3�>.�r�>]��Tݫs�o�:��pQ�<3X�$�W����xi��q� met_�M6}ŠUU���[����t��b��[��$B��xfQ�Z뼉n�E��L����SZ��߅[�s<�{��<wc#'2�(v:�uK�%|-&�C5X
�F�k�-Q�r����EpY.@���[����7��ˣ!�f7�Zo�_S�o�c�{���FvҜ�B��wjz�a��,��0X�Aw*&�C���+fm`s�:�舤���X�Fol�pޘ3Kf����jy�{�g"+R��*'W;2���!�$5h-҇;'k�{��S��_c{x��� v��uޘ�zw<9o6_!���ذqLO��Ѵ��vg��N�Z\{- #������w2�Y�I~�NU�)�D%g'/��B��>�U�W)�P&T�Y�v���#P������:;.�oB{���op�u*.�:=97�kq�ea�A(.�4׍lG�Iʙ�'�"6����;���#ۖAw`���]���ˮ�f�CV�	j-��jBf$e�g����s�������uIm�8�W;��-̳V2�8�q4SK�K(��g �)EKX�0�'�xj� F�3�rv�x��ՀŇuL�B�e�U��'��]�v����&�3qiID������]�`��}y���q;������m��2�_c�\�lꥢՎX��l2��Z�������zz��2�ɐ��^t�s�����{����Y�/g������2�2�V��y��_U��ϻ�]���TiΪ��Y��'�m�A-�ဒf��=�.�����{�V�"���ʦ*0�׹�nM�j��b&hP�G��8j_h�w���.������Q���=����Q��"�.�iEZ{�2>�rF��=؜�.�*�˽U�G��D@�3����'K�hG�Yy���)˹�pb� nѹ�|�ݿ4� !��.0��Z��}K�tuR���]��mK���͔����h�ޝR%�Bn���yTzzJ�h5�*X}�*��R^�A�����+�EY�:��p5�ʛj�R$xw%���6|FƝ�sЙ�������X�$4.�1�ј�����ͨa����V~����e���wC.��j]њ^���C̗��S}���"�	ث1�reH�YpH0KUG|�|�;��o�=W����y+�y�C��E������40`r�=�0�ޡK��l%�ʪ�s�l`�Ӿ<�oʊ��ǋ����j��C��T��"�vmO���cWuM;�uMS��=	{MT�i%��A�X��B�b�w��2 ���K��~�ؽ�����3���{�hUCW;Z���;��}�������SHGGp'�\�Pa"�Wv���Dkʇ��!vK�u��3H�ym_���������'+VA'��K9rٳq�ޥT�5m۾���Q��+(Acy(3W��-��,��6�'�n�,��"�\X����"7�/��Tn&O��ɘ�I����&R�z���&��F2�*�p���^o��n�V���U��Y��n��a#0�ܪ	��\yύUB�M/<|�����ڿ)�~�zz"�e)�I{��WQl���z�zi��3}N�E�誤"3N=}|Y��=��mM.���F<m�`b�v;5Ǆ PZ�!�n	e��@(M����5˺��^�A�C�^7��o>����i��wJ��驈��U�q=V.��xѪ}9ҪR�x����-�`��w����P\��M�1;Y�UE��d磌��9�F/�:�p��h�X�ɔ-M#��?*�f2{Ԅ�0o6�u�*%��#zk&(���x�7ɽ��k���n�zn�1Ц^[�R)�UX�s�n*V]�w�=?�UHҔO�v�dF��ܢp	������^��<�0�X�d���vT��L���,���i��ѿ����ˍ�7��0���TR���Qtn��}|�ߟ�����F�k��n`J�
��m1�G�,ԛ&hD$�ҭG{����'V���J�ھ�8# �/�P�;=��!�����8c�ј��I�����ɵ�(u�٧�Ge�w���TUz	�=�2�'��&oy͋��G����.����ɚ�W��}�R)6Q��8	����E�r�%˺�{�bgݙJ�
̀7��y��<�4B-�!�J�W����$�Љ=1���7j��$�|�is핆���=I,P���	�r�τA�ɘ���&Lթ���`�G�_��V�ƛ+��u���b�)-�]n���[p��-D6˂�?"v;6����7��$�7���`h��D��Z�[�,��]�صs�q�;���H0tu�u'����d��j�ojg#�6X�%��K:�%�m��;\!�wC�S�,�*��M*M���'.�X���u;&zy���d��\��gV�K@���$m�R�ib��Jm/ZO��z�`3�׭C�D�Z<��H�1۶�b�Iѭ�bXKG�#	oN�) R
�h��W�ܖ��t�kֵmϩ�ǘ�s�g������e
�W�{ܪ�5��^�ps�S���B�F�]��ڳ����Ap�Nl�Z�~�>W��;�����!K�m*�
�ʺL!Q+gE��w�$�A8����7 {��,��k����H�>��IwmEm/.��	B�j�%H�n���d�x���0��bS���R��U�b�U5W�δ���ބ�$C�	՛>�𪤍F����<���JKz�@>������)(Y�^wn#:g��@�R���ˋm�3�.�yn��}���+3�;�=���f��d�vtŹ���/{���QS�4!oHI^��h����y=�~���y��~{t�0z�H��8Y�~�.u�d%�h��NW^1囜3Wk��ȶ�z�����׼�p��'3iN��jyZ;u�B RTe�0k�D?�a5c�쯞�e�	j5?}�yӫǢ��.yܭ^���.�dq$�a�hBi��͔=ޚ�U������d�_]�T���3�{�=6�!�pap���"�19]�Yy�>��,��w}5ԅ��r�\Ә�^��i��-�a#UigyUR1*X�{s���u�;�^��c���W�"���P�	��=�h��b�9��딼scnah�j�Ϸ���ĭ؉fM�5|��}r�,���j�l�8z~ރ�4���PC�/t �@'h�u׷�i�9�!���yT^�{ʻ����Ҩ���\i
c���%CA:�7�g�7t���Vx�b���U�O�5T�c��Ý~7��%�X��UI���_��Ѭ��޳�V��]�Vh���Vr�7�~k�����&��(R
��!P�6k�i[9��q\hy;�J~>Z�u���ո����5���-U���1C֮�{Ʀ���f��{F���0�	�3U7�y��0|J$I(BL�E�=|�R?!B5<U�J��T�BW��W�e�[ڍ�y$I��-ӽ{b3��s�z��I��9��Jn��sɧ��z3[�G�=8��O\�(�tj�,�?� ����T�$w�|�/�%�t(�r��"'q�:�7F���2"��꯬}��� /����0Z-�ٿ���M.}҅FѦ��6\���T▽�G^@06!�I�l����o�+qE�^d�H��t�^τ�Q���~u�i�fyCA�r�˝�NɊ&�P�?1�l|�.Z@��_6����L�2x�da�;�����ƣ"詟D1D�%�E��]U���˦l�9�(J�6��RT�^U
U2j�{}W�]��NW�<}�m����Ե*��yt�-�\iٷ����Ǟ�y��]6��^�M�c�E��Z��^lCMuF�X7b�.J�m�������b��I��M� eN1��UH.�N*�y���^�ˋf�Q�>��y�@)�a�D���}�[�Uƚ��X��I���AI߱Ѧ>������)%՗�|�\1#}�c��RF��Sײ4�7���=�������]E���@.iCh�����^%��"g��)u��	����$d�W��*�[q������S� ���1�5F*>���0����ٵ�.D�@{�O�_�؜�R!3��oLA&��-�6c{z$�Um�ʖF�o]l�@�1f�bv�`:Ϋ�t�?l�hv:�\���q��} ��8�[�quEIa	�X�-I��]F2�q��Fڍܒ��nНuu��*����a�G]���L�-H+�����\�܏e�e�6k]��^:����]i��\�.����s%���6�=�L��Sd5�����X�l�G2Q�8��n��s`���:����'�����Opi�����+�ML%]�0 ��q��`�ÒP֖�G꫾m5 '��	(u��u��74����������mm�c��v뵳etţ겇>�e<�RE/j��Ѧ��nbB��t(,�\�%�P)�uh����0G��d�q=��U;�K:xz��9�4=W���0b���A�f�R�V,�>��b�wTzb�㏀=��Lf��gw؋D��S���F�h�iBp�uf�1gn��T(�7���){��֣c���ۂ4��K|<���@d �.*�{g�5v��}фd_�="5_�����x�ڧ��� ���PP�m�AA�̫�m�:�Ch���ڻ��J��{;���t��\�?2������$fl��n�<U�.��������"�o�0S�!(f
u�L-�:j�1�E�:�|��P�Q��p��W��[6�y@6�Zl�����۷�%�������	n����BS������_��X)u�42Tq�)��gșlr���j���f��ڗZ�eխA}� B� @F)W��:�c�����t����;��u���H5
wSf!or����*]���}R戤`_l�3Z�Į$����h^�}ː�v �VTT�L�>֨�Η8[�h5��JO��e����0j��=�?R(}�"V���R��q����QSQ��6g������8�5�(�6�۪��c�W�K.g����3<�_���I���FMJRش��k��m�r�/�^���otl1\�TT�=�0��X�B�]aK=�*��{�d-ۇT�gJ�(,�MVhHFHN=��4���)]�Z{�WG��+!ӡ�#ՠ3˱W�Vy[�i�0V:��j�A:Ԧ�v��UwH�N�pk������_�e�+L�Ly5�*xN�\��g�����5�b�#��kŇ�m��2͍�Y�Px����l�m��r���q�o���.���W��>���:�S��\��3���]�<&kg�`�T���,��Dj�]8��i���e�x" 
9�AsE�RF���p�̀]��z�]9��_<��mr�3���W_R9��ջ�Ͻ�u�;��OQ
�U4Ĩ�,�
�1�����B��=3���_0��`S�O�Y������o�r3V��Uʝa �(wVL�y��Ƽ��z�FX�}�݈�s37Ub~���]�%���4���,�Z��Yo�v��غԸH�댽i���#��Ga���n�v�O�|��=�շ�B�jw�����Vm��������TI���:�$�{3��nL�7�C3;�Z*;cd��]<mz۫���i�S������+\���2L7@GT�^w_bIb����.f�J�
(��4�?W{B8�z陬җ}����]����\���-�
6���Y�#r��`�u
�/&G&�(�a������t�V؅�ja�������4�����㷘����W��6j���l++{�}3�ɳ˻�i��t#/d�s]a��0B�! �/%3Ot3B4U�w`<��e��P���:�Op�ˡQ������ݺL�E}W5���D��ʻ�IrQˍӼ�mWrt]y�{ٹu���h���C��"E[����r��z�V-�.Pё��I�8=�SV���e�R�q^�=�t=}��ʞ�[��L�Ow4}j�����:wM��jb.W�Α�8�hx0���7�"�]��׬x�7�x��|�h�)�>��\�x��T�xo:��8���:!ь�����YyP*\#xo7��`	-<<m������j�~RW�Y�f���zp�Hh��W�jؔF|1�E�g�Yf姵�h�������e�;�-�/f����4�)�7c,@�J�L�b�ٕ��t��w^���p�㹎)��0�AD�A9�Sgi�[guؽ��׉l��,�,��I�����̋��Mej�b�D:��mܮ�c��qۊ�1V���U���[��u�n��)sA�����!��L���o�=N��QX3zk���mS0[Գ�{s2׋��ފ�����k`�bicK@,!N�,��p%O(�N������;����=�ǔ�$���b9���ۗ�ufI��)�F�ƒ� 'N$O���2up!���F�n,� ���JH�W�扡���Tb�9uB�ܽ��6���@d�[-���>�=@���yb.τ�!sS�
��WƐ��	WϷ߿@W�li2p�jq��t�����j8�`��l���-�`�	$� 4�
���Tu^j���]]p�m,����y�Ai�hк�	n�Up�bLu-�!j޼��=�G#֫�^�UgqIC*ǏkE��	�CM�E��Jh+͙���wA�xL��fyO�����)�Q!��ڤmGa�p���N��������]�s�͟Q#�5~��:�7#�&��<S1�S�D`Y*$E��]�Q�?8�,�|�ll<�+rc}J2ک��aU\���'q�V*���-p�2���� 8e�W�q�ǢւZ��N�M\�ʋ��)(�h�v�^z�*�M��댥��=�ϱ��t"h�xD���m���7.�����Nb�vg��z�!g�>�#��0fC�4TYp�4`�i,�+��^7v�{_�~TV����k0�#e��uE���Ȣ��@-R���׳�1xb����τ]�>٦hD,�UT�=�+�mȐ>lz-��o� ��uH�Ǣg݁٠�Ԯ�t�\�tz � �|��+*��^L?E�����{���^��(DH6!d�H�r��'� :H�, �֖w�ɻ�L�؄�>ΗF�g)�F�j�8G�횕Z(`��ӡO
��+�{_�+����S�YN}<h�a��Ʌ��&��sps�td�QL�r>	߼���t32�p� ���c�x���Wm�y4�u���řÇ�>{/�ն�lr�m�]�BM�)���k`(����b|KP�G�F�8����yL]c���"�u��@���Uk�F���.�$�k�#%���y,�u��y���,e�n��jWK]l�I�����&�#rEۀ�l aPC�3�D��$�l)_Pn�I�����W�{d�����[�X`A�\0��e��n��;z�jL�pRJs׶�Q�r�/gnG)C��`2Snk�ϟ��r����To��O���b�+�*�B�vĕ,"ZR�ɵq�鬬`��o'�qMR�ܮ������1�B�E���#� ���b��𛥌>S��"KIyX�ng��^��UB�=�C(%�\U���{çr�{�[���yzz%}�����3�1rkc���|>�ݠ����	4�/<Rɋj��ܘ�վ��V-�|'�������F���ٓhBˊ�����:�tb�h�ce�&��nl�B}m��	p.LQ}��!���m��QTifydБ�o�nb�juӤ���*a$�a2V��(����G����VY$��5�_r�>F�#E	��C}�itN�������jy��q9��F���r�|�׻Ͳ9;jd�~��G'�kyv)�*����r����1cC�~D7�j��_TY��V�|��v�����BE���D����y���'d�s:2��Ա{��7�mC��P��>i�2�I�n��P�?;q�g��s���w�6�y���[��☙5�#�y A,`�M����J���{ܪ6����u�a�?_��W�?=i��F�<eѤ��	���r^j�nŶ�r�+z�h(��/n_�ռs>�=�[�d5F�=ꊣW�P�Rǯʢ'֩R	5��Y�'�_o��<QH ��/�f}�b�c�TY˸�oW���[�?ep��CB�"1��x�-"�!��qu%��1'�\�fxRD����_c����3��R�<���.��!�J�DT
N�gn�a�ztC���h��B^�е'���/+�}Я�[���V����g�&u��5�rc�Ū��Dr0:�t�Hʣj��v�;/*J����C��,������wdW<�S�{�b�W��OP����vi(� ��
0�J*��{�QSHŎ'�>NX��W�������Dt���g͔���-!q�x:3�wv�E�Y�[A�[J}}�ƙ�a(MJ!�M�վ�QF�oV�j���WЈ�� Y��ժ��o�>AB脡A���Xq&;gٵ�a�:�ң{�UK�v�]�8HӚjb�I�o���e�K���W*����?L��[�v��ݘY��P�*[��8m	��)�9�n��Tr9����*��w��	�)�5b<��G�!]E�\BpL=qX�8^�Z�A=0�\vOémdk���ғ��g�8Pg&��)���,T
5(�"%�=�	��R��0�L���U�q�u�@H�p��L|�%���4g��(d�U�W�W�s#������N:1J�]E�>&�b&1����x��n��z���7T�Ǩm�Q��n�޹aߏ�a�AI��6!Vڞ�f
�X���5X����1`�Ꭓuhw>+� LM�wJ�~ޫ� �Ղ����8�7�G��FȏY�W��/��}h�H ��Ž�3�=���bG���g��J�gzf(ҋ�=4�pS��n�:��Y�0�"�_�z��#7� Q�[']���1�?dNR9��$�� i@3WkO�J�������H�t=�F���UP�z����lF������;$P�j���J�E��pF3s��SCsjn[ta����H@{a�mo��,��*^Q��gv��\�6W��ݙ�m=�
;R�����n�a-8��Q��a퍌�����h��U��72g8v�x�\�sZ{mՋ�����k{t����Y�78�z��kC0��3�f٦�ə�1�I����%�8wi�5�W���&�3�9!z�dàqp�7V)bEx�lݝ����PB��瘐��:.E=BX�yF�~<Ni�D�k�`ٸ"L���_I�����aA�Z\��h���c]O\ܻWtv�sN�]Gg�ozN�˗p����{��ER��TP����v���!r�U:KW���!2�9�=�S��8FyI���*�V�7����W{.�8�$����w����l�Y!oOx��?r��M�S~�T[%����.���R��	`8@g���ܦ�}(�r�y%��k��5������Z����MAp�H��4o7�RDQ;~�Gѻ�%7���w�12}�d�0�����H�W5a0�J�Il�0���X��]Q.c6��%�F��`3$�g�\�ު�;�8����mu�[��T>��8�6!W\ݫvc���)���
f��]��5WI[@��t0Fn�B�_e +��V@��ne�ƌ�`�D�ʑBָ����G��_r�]�n>����==0y`2cG�x�+�錍�.h5ę]ƅ��S�{�ے*-g�:�鉨�A���d_
�nE����;��/%\��&�AZ)c��jo~���C;��:�]D{GJ��n��²��kO��'{TUR�;��_�B++�����[ފ��l$�V.�^��ΥLM>6*�{��j,Xk_�Ƞ${E}�K�&V8�pl�$s̉r��"4�Y��;�5�������;ơP�P@N*�!z{��;�uF��?�>B��(�k|f��\��I��@ 0�./0���Q
tGqU�]j�%Z}�QTo^��s���^�$ո%����]�s����]Q�A� O�"�m�s1���4B�1�틅rvcg>N�"Y�:!�(���bv�Kt`������uޠ�FN�T(�KBu��Uy|�qX�Wv�Y޺bc��Q0��M oн4*h.���vͱ�9���&@*�Yk���t]����]�cr��*׼����D�o>���dw�(�(��L�٪=����G���DC-p��U�[�U�:*i��7ǈP��N닳�0^�XH� b��gN�w�>���� ��!�-&�]���qIFs�J�{��m��o�����U�9?OJ*ʵh�m�VR9��#�e����5�����\���7�E�~�Cp�p�,��egr���Gq�܈�jro^?+TWc�Z��sx$�(���_f��"�,y~��i���+�sF�6�D�}���쟬G��]�N��Q0��v�\>��ޫ�cLĞe�X������a�D<_�;�ښ���ҫ�������(1���Va�PJƅ�㢞��N�^�`ט	6`2IB��!���N�tEnw���ߗ�ݘO�zܜL۩��<���D�]�uljn&�����O)��G0���y�-�-��"�I���"2�U��MQAnr�T�_���G���٬�4�Ao�(���P�j.]ߺ|*%������c��Sc0�����١��@��� W�|l&�-S
f�k�3T�e�>���*A3�u�j*�*���B��-5�&����Lz���~t{�T���8L:޻b)#��5G�D�2����K���GW������T�^�+j������#�Q�����#�1��F~��SOq��
⪪��7��0ٙ�N��������8�ܹUw���:�������t[������]L�7�Ǩ��K�����F3H��&͍&m��gccI�4�m�q��7�C��᱙@3��(㎮n8�r�d��fl6t�gUϗ0��mM�f+�F�ے�Fͺ~}ώZ�l6͹t�c3��c���3;3l.\6�m����-�ն��ٸ~��a�f��G0so=ϧ.V;g�ø��<T@pc���`9��@ܑ��D��3Ԩ�{�ٌՍ���V�%[x��(x�r98�:�y�?��+���z���������B���=ῇ��q�zn7o���{ǿ�n���g�v+����EY����x��>#��}_���鿁u�゗�8�<��'�=����p�u�7ё����gX����ί,��|}=�;�yo��\����<'�m�37��M���O���������ߗm�Vr��m�xنo{u�b�l��7�艫6�6���xx��p�|-�]A�m�o�u��9�����ѿ�<����ros|���ӻ�c�S���_6c�lٙ���c���\��������iG�;�����m���B��������ɶ�;ۙa<�����[�qg=��z>#��~v��񣃃��Ӟ~^~=����^��q͜йr��x�\:�����a�>]�g��z9��|[��z7G,�-�g(��$�a�^��G�?�c!���\l�PL\�P���b�Y"l�Yh�P�H��Y�Y[u�pᬋYE��Ɖd��Y��F�(��-4�Ţ�[Ke4m++�d�e�VQL��kl����bֵ����K��(L,Z��E2�-�+$Z%�VZ�4Z�+"-2D�D��E�-de��k,�D�+SQY"�Mk�H�D�QYX�h��Z�H�ZśYEe�"X��Dmd�Eid���6��E4�Ț(�VF�%�%�(�5�+(�B�"l�h�b�+Ye�E��k��VM��"$Ke2Z�Y���Yh�k%�&е�e��$KF��X��,�Y!m�X�D�E	d�lBYYh��"�Q6����E��Ŷ�-��Z+%�,�$�$H�(��m�F�Q,�h�FD��2"�VY�E�E�,�"YEe�����b�,��E4��(Z$[4�BX�F����H���ZMm�Z(�H�Q�̲D��-eV&Ȭ�ڋYEehh���DQk-ȋl�5�VH�H�,Ȣ�E�-�4KZ�d�%�$�E��։b,CE�ZXZ�$[2kE��K-e���VZ%�e�LY"�ĉ��E�e����Ke�Ee�h��E���+$H�V�,ȓQEd��Ɉ���-jɴH�+(��[h�-d���Z%���%��Zb�!&�,�X���j+-b�D�e�,Z%�Z)��b�b��"�-��j-%���LQYB�XX�DQ,��[$Z̢��P�+V%��d$�VQBB��f�&�E	�b"�Z��$QX��Qm�j�+(S-�Yh��Ų+$K�e2̛Q,VH�k-�Q"�Y!,����[kD�,Y��%�VQ,��P�ef����d��5d��P�QL�[Z�j�b4SjQF��Y���&,Z(����$ZX�$K(���M�YX��4&�Sj�e�6��ZĊ-�(�Hk5�j+$K4k-m,�B�6�m�j�f��+(�P���f��,���Z+%�Ų��PQab�B��Dk$Km��[,�Մ���+�kE-�VS(VQ!f��m�k�I�MfE
Ţ�D�6��ebMm��(��++QYX[,���YFDY���VQ,H�YE��QX���V����5�̑EehkX����&��VV��YEb���f�(��6��V�l�V+4���(�(�5f����څ5k$5b�F�aE6�رD�VP���$Kl�aYM��(�VKH�H���%�K%�bDk+4�M��5��EemX�eVQYhP�4������ebE�P���+$-2Y"ū(�S++5�
(��,��"�4�m�
+5b�ɑX�EbM,B�(Vj��++ieVH��Y�-��e����(��d,ZeP����E6��B�"���YdQY,Q"Y��kXSVV��h(V%�"X��VP�M�L��Mej+-f�Qf���+4�[[jSj&�̬�kD�Y�e��+6��$Zm-FB(�V(��6���QmE����YEbEe���Y"����4,V(V%�hQYMEe�D�(�$K!m,���$Zd�b�k5kD�$B�V�-�K(�k+�(�L�k5eڱ�Vi%�Mm�$V%��&��,�X�V�YEjɖj�(X�(ձ!bĲ�&�-�&HVQ,�E��KH���,$K(��em,��h�K!m�QY"�S+VYlՖ�d"��[��ji�d�fH��)�9x�1ɵl։�QH�P�D�Qk(���,V)�Z�+��l��bXVB$QEef�VM6S(���h�VHV%�Ȗej(�4ڍEb���(�h�[)��e��(�++	+$VS5�+5�h��+(��Ee�+(���mMh�Ք+4E6Qk$V��2�E3[",Պ+([XQ[d#VQY�(��
�,Qm1B,��AM�4,�I�b"���m,���°�Y���
-b�V����j-���(в���,Z%�Ed��$)���$V(��QB�Eef��LQYf�D�E2�md$-b���JZ�ҍE%X��%��%UV6ԫ[T�&���R�*RkU�mIJJV�k)U&����R�E�UI*[%,��L��6�դ�U���I���T�J[U���$��Je�Q*��Md��%"�B*���VԫMUU�J��B�,������%e�3eUV�V��D���V�U���J�*�lZ�ԒZ���+-5J�T�EZ�) �$ҥV�)�Jҥ+*�YKYZ�d�UeRDT�U��mR��T�mR�A���nI����ke����e�VҖe�T���ij�J�UJ�JVDJ�ғm��k*���-+YU-b��U*�UJ�m�����Z�SUR���CeZ�*"�j�Ȳʚ�)jZ���k[YdZ������V�E�����"J�TYY�m�ȷM[��Q*�-+"Z�J[J�6UUT�"�kRJ�*�e�%kl�T�KYkKT��Z�"E�e����,�5�E�eDU���Ie*�*ֲ�m��V�Z�K$L�J��j�U�i��ҵ$�b+R�Y"��(�d��*DYT���j�6md��Z���)��EY�Z�VH���������"%j,���VQJFڭe�k-���Z3Mh�ZR�Ȋ�!6Ȭ��EdEe6����"QD�V�3YkDVKT�JH����Vֲ-R"*�DFMMK"�Qh�Q6֫,�e�Z-
*-E&d��EV։�*���dl�dE�VKY�E��dJ�d�*ZD���#4-(�U�ZY��Q,��K(��E��J�(��Z��YD�d�Yh�"�3,��Q[UK�l�D�"�d�Y[��a�%�K+iee�dص��,�$QME�Ee�%�mՒ+(�Yh��D�m",Ye��+%���[(��X�(�15�DZ�Qh�C,�h�-$H�Z,Œ%��ښ��-���h�E26�d�e��-Y)�QY"X[bŢ�e�,��Yf�D��e��-�Z+�Q,�V�X�H���F�h�Q,�YE5�Z+$VQEe�6�-,ֲ�m�'Ι���Zi UATh���H��&(,����0�3r���w�7�z���Mѿ�f���m�n�9��;z�O�M�o��|����<6���;w��|��ltÓq�Q�oGk:��޷�&���-��=���u�ն�GMٛy��t[�`<������ߓl��w���ݽ��~��27�r��3uF8�q�m�������͞�ǳ��p��s�~?���w7F�}[�n���6�]{���n͟��}=��M�i�Q3�<������z8���g�u�gwɿ3�nǩ��6ٙ��'�;�ͳՋ4˖<[�`�ɾ��bO����ξ��s�'+u�w��>m�!�[&��ۺz�m�ٙ��K��f�����|���[okk}G_߬�k���m�r:f�:7���n��_Gsv���6�n���3�����3u��f�Ǵ��8kM�aͫ\nc���6��iϵ8&�l�fY��n�w��=��6�ϓ�m�v��ۗ#�-����9�3�ۍ��3�g���7�v��ݞ%�V�έ���	bA#3�:��9I���;�$C�v����l��nC�ޛ���>A�xl/����;[߳ffo��o�����O~v{1�ͨ����^�<�[�gǾ�7��x��?����9���3�oI����O-�c��V�Ǐ��un1o��C��ܾm��kr���om�7ɿ1Λ�5��u��ocͷ��ߺ�����͙��9���>Vz~#����X����:�ˎ�X��ٙ��ێA��G�#�[��'w6ތ�|�yQ��3�z6n�-�vׇv��n۵�[#�,���Я��I�� �QD�D��?��7Ǻ������̶Qr�7o���;��#B&�|�};�|��c���n�,�.8N:ov��9�畭��7W������ٳ34y[���[��=L��|.5��Y�;7�z�����n7�n��6�|�}����ַ��z6�;�c:k|��E�'�pܹ^��t[���p�޳���-�na��G1/W}y�n�t�w�m��g�{C���7����oǩ�f����ۡ���m�iS�u�^wtOK�30�����;�=�y�7Woft��q�]��X����u�r�\��·_l�Q՟�������S�8᳞F���"m������{����H�
�>�`